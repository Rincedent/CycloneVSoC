-- standalone_hps.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity standalone_hps is
	port (
		buttons_i_export                : in    std_logic_vector(3 downto 0)  := (others => '0'); -- buttons_i.export
		clk_clk                         : in    std_logic                     := '0';             --       clk.clk
		dipsw_i_export                  : in    std_logic_vector(3 downto 0)  := (others => '0'); --   dipsw_i.export
		h2f_bus_awid                    : out   std_logic_vector(11 downto 0);                    --   h2f_bus.awid
		h2f_bus_awaddr                  : out   std_logic_vector(29 downto 0);                    --          .awaddr
		h2f_bus_awlen                   : out   std_logic_vector(7 downto 0);                     --          .awlen
		h2f_bus_awsize                  : out   std_logic_vector(2 downto 0);                     --          .awsize
		h2f_bus_awburst                 : out   std_logic_vector(1 downto 0);                     --          .awburst
		h2f_bus_awlock                  : out   std_logic_vector(0 downto 0);                     --          .awlock
		h2f_bus_awcache                 : out   std_logic_vector(3 downto 0);                     --          .awcache
		h2f_bus_awprot                  : out   std_logic_vector(2 downto 0);                     --          .awprot
		h2f_bus_awqos                   : out   std_logic_vector(3 downto 0);                     --          .awqos
		h2f_bus_awvalid                 : out   std_logic;                                        --          .awvalid
		h2f_bus_awready                 : in    std_logic                     := '0';             --          .awready
		h2f_bus_wdata                   : out   std_logic_vector(31 downto 0);                    --          .wdata
		h2f_bus_wstrb                   : out   std_logic_vector(3 downto 0);                     --          .wstrb
		h2f_bus_wlast                   : out   std_logic;                                        --          .wlast
		h2f_bus_wvalid                  : out   std_logic;                                        --          .wvalid
		h2f_bus_wready                  : in    std_logic                     := '0';             --          .wready
		h2f_bus_bid                     : in    std_logic_vector(11 downto 0) := (others => '0'); --          .bid
		h2f_bus_bresp                   : in    std_logic_vector(1 downto 0)  := (others => '0'); --          .bresp
		h2f_bus_bvalid                  : in    std_logic                     := '0';             --          .bvalid
		h2f_bus_bready                  : out   std_logic;                                        --          .bready
		h2f_bus_arid                    : out   std_logic_vector(11 downto 0);                    --          .arid
		h2f_bus_araddr                  : out   std_logic_vector(29 downto 0);                    --          .araddr
		h2f_bus_arlen                   : out   std_logic_vector(7 downto 0);                     --          .arlen
		h2f_bus_arsize                  : out   std_logic_vector(2 downto 0);                     --          .arsize
		h2f_bus_arburst                 : out   std_logic_vector(1 downto 0);                     --          .arburst
		h2f_bus_arlock                  : out   std_logic_vector(0 downto 0);                     --          .arlock
		h2f_bus_arcache                 : out   std_logic_vector(3 downto 0);                     --          .arcache
		h2f_bus_arprot                  : out   std_logic_vector(2 downto 0);                     --          .arprot
		h2f_bus_arqos                   : out   std_logic_vector(3 downto 0);                     --          .arqos
		h2f_bus_arvalid                 : out   std_logic;                                        --          .arvalid
		h2f_bus_arready                 : in    std_logic                     := '0';             --          .arready
		h2f_bus_rid                     : in    std_logic_vector(11 downto 0) := (others => '0'); --          .rid
		h2f_bus_rdata                   : in    std_logic_vector(31 downto 0) := (others => '0'); --          .rdata
		h2f_bus_rresp                   : in    std_logic_vector(1 downto 0)  := (others => '0'); --          .rresp
		h2f_bus_rlast                   : in    std_logic                     := '0';             --          .rlast
		h2f_bus_rvalid                  : in    std_logic                     := '0';             --          .rvalid
		h2f_bus_rready                  : out   std_logic;                                        --          .rready
		h2f_reset_reset_n               : out   std_logic;                                        -- h2f_reset.reset_n
		hps_io_hps_io_emac1_inst_TX_CLK : out   std_logic;                                        --    hps_io.hps_io_emac1_inst_TX_CLK
		hps_io_hps_io_emac1_inst_TXD0   : out   std_logic;                                        --          .hps_io_emac1_inst_TXD0
		hps_io_hps_io_emac1_inst_TXD1   : out   std_logic;                                        --          .hps_io_emac1_inst_TXD1
		hps_io_hps_io_emac1_inst_TXD2   : out   std_logic;                                        --          .hps_io_emac1_inst_TXD2
		hps_io_hps_io_emac1_inst_TXD3   : out   std_logic;                                        --          .hps_io_emac1_inst_TXD3
		hps_io_hps_io_emac1_inst_RXD0   : in    std_logic                     := '0';             --          .hps_io_emac1_inst_RXD0
		hps_io_hps_io_emac1_inst_MDIO   : inout std_logic                     := '0';             --          .hps_io_emac1_inst_MDIO
		hps_io_hps_io_emac1_inst_MDC    : out   std_logic;                                        --          .hps_io_emac1_inst_MDC
		hps_io_hps_io_emac1_inst_RX_CTL : in    std_logic                     := '0';             --          .hps_io_emac1_inst_RX_CTL
		hps_io_hps_io_emac1_inst_TX_CTL : out   std_logic;                                        --          .hps_io_emac1_inst_TX_CTL
		hps_io_hps_io_emac1_inst_RX_CLK : in    std_logic                     := '0';             --          .hps_io_emac1_inst_RX_CLK
		hps_io_hps_io_emac1_inst_RXD1   : in    std_logic                     := '0';             --          .hps_io_emac1_inst_RXD1
		hps_io_hps_io_emac1_inst_RXD2   : in    std_logic                     := '0';             --          .hps_io_emac1_inst_RXD2
		hps_io_hps_io_emac1_inst_RXD3   : in    std_logic                     := '0';             --          .hps_io_emac1_inst_RXD3
		hps_io_hps_io_qspi_inst_IO0     : inout std_logic                     := '0';             --          .hps_io_qspi_inst_IO0
		hps_io_hps_io_qspi_inst_IO1     : inout std_logic                     := '0';             --          .hps_io_qspi_inst_IO1
		hps_io_hps_io_qspi_inst_IO2     : inout std_logic                     := '0';             --          .hps_io_qspi_inst_IO2
		hps_io_hps_io_qspi_inst_IO3     : inout std_logic                     := '0';             --          .hps_io_qspi_inst_IO3
		hps_io_hps_io_qspi_inst_SS0     : out   std_logic;                                        --          .hps_io_qspi_inst_SS0
		hps_io_hps_io_qspi_inst_CLK     : out   std_logic;                                        --          .hps_io_qspi_inst_CLK
		hps_io_hps_io_sdio_inst_CMD     : inout std_logic                     := '0';             --          .hps_io_sdio_inst_CMD
		hps_io_hps_io_sdio_inst_D0      : inout std_logic                     := '0';             --          .hps_io_sdio_inst_D0
		hps_io_hps_io_sdio_inst_D1      : inout std_logic                     := '0';             --          .hps_io_sdio_inst_D1
		hps_io_hps_io_sdio_inst_CLK     : out   std_logic;                                        --          .hps_io_sdio_inst_CLK
		hps_io_hps_io_sdio_inst_D2      : inout std_logic                     := '0';             --          .hps_io_sdio_inst_D2
		hps_io_hps_io_sdio_inst_D3      : inout std_logic                     := '0';             --          .hps_io_sdio_inst_D3
		hps_io_hps_io_usb1_inst_D0      : inout std_logic                     := '0';             --          .hps_io_usb1_inst_D0
		hps_io_hps_io_usb1_inst_D1      : inout std_logic                     := '0';             --          .hps_io_usb1_inst_D1
		hps_io_hps_io_usb1_inst_D2      : inout std_logic                     := '0';             --          .hps_io_usb1_inst_D2
		hps_io_hps_io_usb1_inst_D3      : inout std_logic                     := '0';             --          .hps_io_usb1_inst_D3
		hps_io_hps_io_usb1_inst_D4      : inout std_logic                     := '0';             --          .hps_io_usb1_inst_D4
		hps_io_hps_io_usb1_inst_D5      : inout std_logic                     := '0';             --          .hps_io_usb1_inst_D5
		hps_io_hps_io_usb1_inst_D6      : inout std_logic                     := '0';             --          .hps_io_usb1_inst_D6
		hps_io_hps_io_usb1_inst_D7      : inout std_logic                     := '0';             --          .hps_io_usb1_inst_D7
		hps_io_hps_io_usb1_inst_CLK     : in    std_logic                     := '0';             --          .hps_io_usb1_inst_CLK
		hps_io_hps_io_usb1_inst_STP     : out   std_logic;                                        --          .hps_io_usb1_inst_STP
		hps_io_hps_io_usb1_inst_DIR     : in    std_logic                     := '0';             --          .hps_io_usb1_inst_DIR
		hps_io_hps_io_usb1_inst_NXT     : in    std_logic                     := '0';             --          .hps_io_usb1_inst_NXT
		hps_io_hps_io_spim0_inst_CLK    : out   std_logic;                                        --          .hps_io_spim0_inst_CLK
		hps_io_hps_io_spim0_inst_MOSI   : out   std_logic;                                        --          .hps_io_spim0_inst_MOSI
		hps_io_hps_io_spim0_inst_MISO   : in    std_logic                     := '0';             --          .hps_io_spim0_inst_MISO
		hps_io_hps_io_spim0_inst_SS0    : out   std_logic;                                        --          .hps_io_spim0_inst_SS0
		hps_io_hps_io_uart0_inst_RX     : in    std_logic                     := '0';             --          .hps_io_uart0_inst_RX
		hps_io_hps_io_uart0_inst_TX     : out   std_logic;                                        --          .hps_io_uart0_inst_TX
		hps_io_hps_io_i2c0_inst_SDA     : inout std_logic                     := '0';             --          .hps_io_i2c0_inst_SDA
		hps_io_hps_io_i2c0_inst_SCL     : inout std_logic                     := '0';             --          .hps_io_i2c0_inst_SCL
		hps_io_hps_io_can0_inst_RX      : in    std_logic                     := '0';             --          .hps_io_can0_inst_RX
		hps_io_hps_io_can0_inst_TX      : out   std_logic;                                        --          .hps_io_can0_inst_TX
		hps_io_hps_io_trace_inst_CLK    : out   std_logic;                                        --          .hps_io_trace_inst_CLK
		hps_io_hps_io_trace_inst_D0     : out   std_logic;                                        --          .hps_io_trace_inst_D0
		hps_io_hps_io_trace_inst_D1     : out   std_logic;                                        --          .hps_io_trace_inst_D1
		hps_io_hps_io_trace_inst_D2     : out   std_logic;                                        --          .hps_io_trace_inst_D2
		hps_io_hps_io_trace_inst_D3     : out   std_logic;                                        --          .hps_io_trace_inst_D3
		hps_io_hps_io_trace_inst_D4     : out   std_logic;                                        --          .hps_io_trace_inst_D4
		hps_io_hps_io_trace_inst_D5     : out   std_logic;                                        --          .hps_io_trace_inst_D5
		hps_io_hps_io_trace_inst_D6     : out   std_logic;                                        --          .hps_io_trace_inst_D6
		hps_io_hps_io_trace_inst_D7     : out   std_logic;                                        --          .hps_io_trace_inst_D7
		leds_o_export                   : out   std_logic_vector(3 downto 0);                     --    leds_o.export
		memory_mem_a                    : out   std_logic_vector(14 downto 0);                    --    memory.mem_a
		memory_mem_ba                   : out   std_logic_vector(2 downto 0);                     --          .mem_ba
		memory_mem_ck                   : out   std_logic;                                        --          .mem_ck
		memory_mem_ck_n                 : out   std_logic;                                        --          .mem_ck_n
		memory_mem_cke                  : out   std_logic;                                        --          .mem_cke
		memory_mem_cs_n                 : out   std_logic;                                        --          .mem_cs_n
		memory_mem_ras_n                : out   std_logic;                                        --          .mem_ras_n
		memory_mem_cas_n                : out   std_logic;                                        --          .mem_cas_n
		memory_mem_we_n                 : out   std_logic;                                        --          .mem_we_n
		memory_mem_reset_n              : out   std_logic;                                        --          .mem_reset_n
		memory_mem_dq                   : inout std_logic_vector(39 downto 0) := (others => '0'); --          .mem_dq
		memory_mem_dqs                  : inout std_logic_vector(4 downto 0)  := (others => '0'); --          .mem_dqs
		memory_mem_dqs_n                : inout std_logic_vector(4 downto 0)  := (others => '0'); --          .mem_dqs_n
		memory_mem_odt                  : out   std_logic;                                        --          .mem_odt
		memory_mem_dm                   : out   std_logic_vector(4 downto 0);                     --          .mem_dm
		memory_oct_rzqin                : in    std_logic                     := '0';             --          .oct_rzqin
		reset_reset_n                   : in    std_logic                     := '0'              --     reset.reset_n
	);
end entity standalone_hps;

architecture rtl of standalone_hps is
	component altera_axi_bridge is
		generic (
			USE_PIPELINE          : integer := 1;
			USE_M0_AWID           : integer := 1;
			USE_M0_AWREGION       : integer := 1;
			USE_M0_AWLEN          : integer := 1;
			USE_M0_AWSIZE         : integer := 1;
			USE_M0_AWBURST        : integer := 1;
			USE_M0_AWLOCK         : integer := 1;
			USE_M0_AWCACHE        : integer := 1;
			USE_M0_AWQOS          : integer := 1;
			USE_S0_AWREGION       : integer := 1;
			USE_S0_AWLOCK         : integer := 1;
			USE_S0_AWCACHE        : integer := 1;
			USE_S0_AWQOS          : integer := 1;
			USE_S0_AWPROT         : integer := 1;
			USE_M0_WSTRB          : integer := 1;
			USE_S0_WLAST          : integer := 1;
			USE_M0_BID            : integer := 1;
			USE_M0_BRESP          : integer := 1;
			USE_S0_BRESP          : integer := 1;
			USE_M0_ARID           : integer := 1;
			USE_M0_ARREGION       : integer := 1;
			USE_M0_ARLEN          : integer := 1;
			USE_M0_ARSIZE         : integer := 1;
			USE_M0_ARBURST        : integer := 1;
			USE_M0_ARLOCK         : integer := 1;
			USE_M0_ARCACHE        : integer := 1;
			USE_M0_ARQOS          : integer := 1;
			USE_S0_ARREGION       : integer := 1;
			USE_S0_ARLOCK         : integer := 1;
			USE_S0_ARCACHE        : integer := 1;
			USE_S0_ARQOS          : integer := 1;
			USE_S0_ARPROT         : integer := 1;
			USE_M0_RID            : integer := 1;
			USE_M0_RRESP          : integer := 1;
			USE_M0_RLAST          : integer := 1;
			USE_S0_RRESP          : integer := 1;
			M0_ID_WIDTH           : integer := 8;
			S0_ID_WIDTH           : integer := 8;
			DATA_WIDTH            : integer := 32;
			WRITE_ADDR_USER_WIDTH : integer := 64;
			READ_ADDR_USER_WIDTH  : integer := 64;
			WRITE_DATA_USER_WIDTH : integer := 64;
			WRITE_RESP_USER_WIDTH : integer := 64;
			READ_DATA_USER_WIDTH  : integer := 64;
			ADDR_WIDTH            : integer := 11;
			USE_S0_AWUSER         : integer := 0;
			USE_S0_ARUSER         : integer := 0;
			USE_S0_WUSER          : integer := 0;
			USE_S0_RUSER          : integer := 0;
			USE_S0_BUSER          : integer := 0;
			USE_M0_AWUSER         : integer := 0;
			USE_M0_ARUSER         : integer := 0;
			USE_M0_WUSER          : integer := 0;
			USE_M0_RUSER          : integer := 0;
			USE_M0_BUSER          : integer := 0;
			AXI_VERSION           : string  := "AXI3";
			BURST_LENGTH_WIDTH    : integer := 4;
			LOCK_WIDTH            : integer := 2
		);
		port (
			aclk        : in  std_logic                     := 'X';             -- clk
			aresetn     : in  std_logic                     := 'X';             -- reset_n
			s0_awid     : in  std_logic_vector(11 downto 0) := (others => 'X'); -- awid
			s0_awaddr   : in  std_logic_vector(29 downto 0) := (others => 'X'); -- awaddr
			s0_awlen    : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- awlen
			s0_awsize   : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- awsize
			s0_awburst  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- awburst
			s0_awlock   : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- awlock
			s0_awcache  : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- awcache
			s0_awprot   : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- awprot
			s0_awqos    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- awqos
			s0_awvalid  : in  std_logic                     := 'X';             -- awvalid
			s0_awready  : out std_logic;                                        -- awready
			s0_wdata    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- wdata
			s0_wstrb    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- wstrb
			s0_wlast    : in  std_logic                     := 'X';             -- wlast
			s0_wvalid   : in  std_logic                     := 'X';             -- wvalid
			s0_wready   : out std_logic;                                        -- wready
			s0_bid      : out std_logic_vector(11 downto 0);                    -- bid
			s0_bresp    : out std_logic_vector(1 downto 0);                     -- bresp
			s0_bvalid   : out std_logic;                                        -- bvalid
			s0_bready   : in  std_logic                     := 'X';             -- bready
			s0_arid     : in  std_logic_vector(11 downto 0) := (others => 'X'); -- arid
			s0_araddr   : in  std_logic_vector(29 downto 0) := (others => 'X'); -- araddr
			s0_arlen    : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- arlen
			s0_arsize   : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- arsize
			s0_arburst  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- arburst
			s0_arlock   : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- arlock
			s0_arcache  : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- arcache
			s0_arprot   : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- arprot
			s0_arqos    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- arqos
			s0_arvalid  : in  std_logic                     := 'X';             -- arvalid
			s0_arready  : out std_logic;                                        -- arready
			s0_rid      : out std_logic_vector(11 downto 0);                    -- rid
			s0_rdata    : out std_logic_vector(31 downto 0);                    -- rdata
			s0_rresp    : out std_logic_vector(1 downto 0);                     -- rresp
			s0_rlast    : out std_logic;                                        -- rlast
			s0_rvalid   : out std_logic;                                        -- rvalid
			s0_rready   : in  std_logic                     := 'X';             -- rready
			m0_awid     : out std_logic_vector(11 downto 0);                    -- awid
			m0_awaddr   : out std_logic_vector(29 downto 0);                    -- awaddr
			m0_awlen    : out std_logic_vector(7 downto 0);                     -- awlen
			m0_awsize   : out std_logic_vector(2 downto 0);                     -- awsize
			m0_awburst  : out std_logic_vector(1 downto 0);                     -- awburst
			m0_awlock   : out std_logic_vector(0 downto 0);                     -- awlock
			m0_awcache  : out std_logic_vector(3 downto 0);                     -- awcache
			m0_awprot   : out std_logic_vector(2 downto 0);                     -- awprot
			m0_awqos    : out std_logic_vector(3 downto 0);                     -- awqos
			m0_awvalid  : out std_logic;                                        -- awvalid
			m0_awready  : in  std_logic                     := 'X';             -- awready
			m0_wdata    : out std_logic_vector(31 downto 0);                    -- wdata
			m0_wstrb    : out std_logic_vector(3 downto 0);                     -- wstrb
			m0_wlast    : out std_logic;                                        -- wlast
			m0_wvalid   : out std_logic;                                        -- wvalid
			m0_wready   : in  std_logic                     := 'X';             -- wready
			m0_bid      : in  std_logic_vector(11 downto 0) := (others => 'X'); -- bid
			m0_bresp    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- bresp
			m0_bvalid   : in  std_logic                     := 'X';             -- bvalid
			m0_bready   : out std_logic;                                        -- bready
			m0_arid     : out std_logic_vector(11 downto 0);                    -- arid
			m0_araddr   : out std_logic_vector(29 downto 0);                    -- araddr
			m0_arlen    : out std_logic_vector(7 downto 0);                     -- arlen
			m0_arsize   : out std_logic_vector(2 downto 0);                     -- arsize
			m0_arburst  : out std_logic_vector(1 downto 0);                     -- arburst
			m0_arlock   : out std_logic_vector(0 downto 0);                     -- arlock
			m0_arcache  : out std_logic_vector(3 downto 0);                     -- arcache
			m0_arprot   : out std_logic_vector(2 downto 0);                     -- arprot
			m0_arqos    : out std_logic_vector(3 downto 0);                     -- arqos
			m0_arvalid  : out std_logic;                                        -- arvalid
			m0_arready  : in  std_logic                     := 'X';             -- arready
			m0_rid      : in  std_logic_vector(11 downto 0) := (others => 'X'); -- rid
			m0_rdata    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- rdata
			m0_rresp    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- rresp
			m0_rlast    : in  std_logic                     := 'X';             -- rlast
			m0_rvalid   : in  std_logic                     := 'X';             -- rvalid
			m0_rready   : out std_logic;                                        -- rready
			s0_awuser   : in  std_logic_vector(63 downto 0) := (others => 'X'); -- awuser
			s0_awregion : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- awregion
			s0_wuser    : in  std_logic_vector(63 downto 0) := (others => 'X'); -- wuser
			s0_buser    : out std_logic_vector(63 downto 0);                    -- buser
			s0_aruser   : in  std_logic_vector(63 downto 0) := (others => 'X'); -- aruser
			s0_arregion : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- arregion
			s0_ruser    : out std_logic_vector(63 downto 0);                    -- ruser
			m0_awuser   : out std_logic_vector(63 downto 0);                    -- awuser
			m0_awregion : out std_logic_vector(3 downto 0);                     -- awregion
			m0_wuser    : out std_logic_vector(63 downto 0);                    -- wuser
			m0_buser    : in  std_logic_vector(63 downto 0) := (others => 'X'); -- buser
			m0_aruser   : out std_logic_vector(63 downto 0);                    -- aruser
			m0_arregion : out std_logic_vector(3 downto 0);                     -- arregion
			m0_ruser    : in  std_logic_vector(63 downto 0) := (others => 'X'); -- ruser
			m0_wid      : out std_logic_vector(11 downto 0);                    -- m0_wid
			s0_wid      : in  std_logic_vector(11 downto 0) := (others => 'X')  -- s0_wid
		);
	end component altera_axi_bridge;

	component standalone_hps_buttons_i is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(3 downto 0)  := (others => 'X')  -- export
		);
	end component standalone_hps_buttons_i;

	component standalone_hps_hps_0 is
		generic (
			F2S_Width : integer := 2;
			S2F_Width : integer := 2
		);
		port (
			f2h_cold_rst_req_n       : in    std_logic                     := 'X';             -- reset_n
			f2h_dbg_rst_req_n        : in    std_logic                     := 'X';             -- reset_n
			f2h_warm_rst_req_n       : in    std_logic                     := 'X';             -- reset_n
			f2h_stm_hwevents         : in    std_logic_vector(27 downto 0) := (others => 'X'); -- stm_hwevents
			mem_a                    : out   std_logic_vector(14 downto 0);                    -- mem_a
			mem_ba                   : out   std_logic_vector(2 downto 0);                     -- mem_ba
			mem_ck                   : out   std_logic;                                        -- mem_ck
			mem_ck_n                 : out   std_logic;                                        -- mem_ck_n
			mem_cke                  : out   std_logic;                                        -- mem_cke
			mem_cs_n                 : out   std_logic;                                        -- mem_cs_n
			mem_ras_n                : out   std_logic;                                        -- mem_ras_n
			mem_cas_n                : out   std_logic;                                        -- mem_cas_n
			mem_we_n                 : out   std_logic;                                        -- mem_we_n
			mem_reset_n              : out   std_logic;                                        -- mem_reset_n
			mem_dq                   : inout std_logic_vector(39 downto 0) := (others => 'X'); -- mem_dq
			mem_dqs                  : inout std_logic_vector(4 downto 0)  := (others => 'X'); -- mem_dqs
			mem_dqs_n                : inout std_logic_vector(4 downto 0)  := (others => 'X'); -- mem_dqs_n
			mem_odt                  : out   std_logic;                                        -- mem_odt
			mem_dm                   : out   std_logic_vector(4 downto 0);                     -- mem_dm
			oct_rzqin                : in    std_logic                     := 'X';             -- oct_rzqin
			hps_io_emac1_inst_TX_CLK : out   std_logic;                                        -- hps_io_emac1_inst_TX_CLK
			hps_io_emac1_inst_TXD0   : out   std_logic;                                        -- hps_io_emac1_inst_TXD0
			hps_io_emac1_inst_TXD1   : out   std_logic;                                        -- hps_io_emac1_inst_TXD1
			hps_io_emac1_inst_TXD2   : out   std_logic;                                        -- hps_io_emac1_inst_TXD2
			hps_io_emac1_inst_TXD3   : out   std_logic;                                        -- hps_io_emac1_inst_TXD3
			hps_io_emac1_inst_RXD0   : in    std_logic                     := 'X';             -- hps_io_emac1_inst_RXD0
			hps_io_emac1_inst_MDIO   : inout std_logic                     := 'X';             -- hps_io_emac1_inst_MDIO
			hps_io_emac1_inst_MDC    : out   std_logic;                                        -- hps_io_emac1_inst_MDC
			hps_io_emac1_inst_RX_CTL : in    std_logic                     := 'X';             -- hps_io_emac1_inst_RX_CTL
			hps_io_emac1_inst_TX_CTL : out   std_logic;                                        -- hps_io_emac1_inst_TX_CTL
			hps_io_emac1_inst_RX_CLK : in    std_logic                     := 'X';             -- hps_io_emac1_inst_RX_CLK
			hps_io_emac1_inst_RXD1   : in    std_logic                     := 'X';             -- hps_io_emac1_inst_RXD1
			hps_io_emac1_inst_RXD2   : in    std_logic                     := 'X';             -- hps_io_emac1_inst_RXD2
			hps_io_emac1_inst_RXD3   : in    std_logic                     := 'X';             -- hps_io_emac1_inst_RXD3
			hps_io_qspi_inst_IO0     : inout std_logic                     := 'X';             -- hps_io_qspi_inst_IO0
			hps_io_qspi_inst_IO1     : inout std_logic                     := 'X';             -- hps_io_qspi_inst_IO1
			hps_io_qspi_inst_IO2     : inout std_logic                     := 'X';             -- hps_io_qspi_inst_IO2
			hps_io_qspi_inst_IO3     : inout std_logic                     := 'X';             -- hps_io_qspi_inst_IO3
			hps_io_qspi_inst_SS0     : out   std_logic;                                        -- hps_io_qspi_inst_SS0
			hps_io_qspi_inst_CLK     : out   std_logic;                                        -- hps_io_qspi_inst_CLK
			hps_io_sdio_inst_CMD     : inout std_logic                     := 'X';             -- hps_io_sdio_inst_CMD
			hps_io_sdio_inst_D0      : inout std_logic                     := 'X';             -- hps_io_sdio_inst_D0
			hps_io_sdio_inst_D1      : inout std_logic                     := 'X';             -- hps_io_sdio_inst_D1
			hps_io_sdio_inst_CLK     : out   std_logic;                                        -- hps_io_sdio_inst_CLK
			hps_io_sdio_inst_D2      : inout std_logic                     := 'X';             -- hps_io_sdio_inst_D2
			hps_io_sdio_inst_D3      : inout std_logic                     := 'X';             -- hps_io_sdio_inst_D3
			hps_io_usb1_inst_D0      : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D0
			hps_io_usb1_inst_D1      : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D1
			hps_io_usb1_inst_D2      : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D2
			hps_io_usb1_inst_D3      : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D3
			hps_io_usb1_inst_D4      : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D4
			hps_io_usb1_inst_D5      : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D5
			hps_io_usb1_inst_D6      : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D6
			hps_io_usb1_inst_D7      : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D7
			hps_io_usb1_inst_CLK     : in    std_logic                     := 'X';             -- hps_io_usb1_inst_CLK
			hps_io_usb1_inst_STP     : out   std_logic;                                        -- hps_io_usb1_inst_STP
			hps_io_usb1_inst_DIR     : in    std_logic                     := 'X';             -- hps_io_usb1_inst_DIR
			hps_io_usb1_inst_NXT     : in    std_logic                     := 'X';             -- hps_io_usb1_inst_NXT
			hps_io_spim0_inst_CLK    : out   std_logic;                                        -- hps_io_spim0_inst_CLK
			hps_io_spim0_inst_MOSI   : out   std_logic;                                        -- hps_io_spim0_inst_MOSI
			hps_io_spim0_inst_MISO   : in    std_logic                     := 'X';             -- hps_io_spim0_inst_MISO
			hps_io_spim0_inst_SS0    : out   std_logic;                                        -- hps_io_spim0_inst_SS0
			hps_io_uart0_inst_RX     : in    std_logic                     := 'X';             -- hps_io_uart0_inst_RX
			hps_io_uart0_inst_TX     : out   std_logic;                                        -- hps_io_uart0_inst_TX
			hps_io_i2c0_inst_SDA     : inout std_logic                     := 'X';             -- hps_io_i2c0_inst_SDA
			hps_io_i2c0_inst_SCL     : inout std_logic                     := 'X';             -- hps_io_i2c0_inst_SCL
			hps_io_can0_inst_RX      : in    std_logic                     := 'X';             -- hps_io_can0_inst_RX
			hps_io_can0_inst_TX      : out   std_logic;                                        -- hps_io_can0_inst_TX
			hps_io_trace_inst_CLK    : out   std_logic;                                        -- hps_io_trace_inst_CLK
			hps_io_trace_inst_D0     : out   std_logic;                                        -- hps_io_trace_inst_D0
			hps_io_trace_inst_D1     : out   std_logic;                                        -- hps_io_trace_inst_D1
			hps_io_trace_inst_D2     : out   std_logic;                                        -- hps_io_trace_inst_D2
			hps_io_trace_inst_D3     : out   std_logic;                                        -- hps_io_trace_inst_D3
			hps_io_trace_inst_D4     : out   std_logic;                                        -- hps_io_trace_inst_D4
			hps_io_trace_inst_D5     : out   std_logic;                                        -- hps_io_trace_inst_D5
			hps_io_trace_inst_D6     : out   std_logic;                                        -- hps_io_trace_inst_D6
			hps_io_trace_inst_D7     : out   std_logic;                                        -- hps_io_trace_inst_D7
			h2f_rst_n                : out   std_logic;                                        -- reset_n
			h2f_axi_clk              : in    std_logic                     := 'X';             -- clk
			h2f_AWID                 : out   std_logic_vector(11 downto 0);                    -- awid
			h2f_AWADDR               : out   std_logic_vector(29 downto 0);                    -- awaddr
			h2f_AWLEN                : out   std_logic_vector(3 downto 0);                     -- awlen
			h2f_AWSIZE               : out   std_logic_vector(2 downto 0);                     -- awsize
			h2f_AWBURST              : out   std_logic_vector(1 downto 0);                     -- awburst
			h2f_AWLOCK               : out   std_logic_vector(1 downto 0);                     -- awlock
			h2f_AWCACHE              : out   std_logic_vector(3 downto 0);                     -- awcache
			h2f_AWPROT               : out   std_logic_vector(2 downto 0);                     -- awprot
			h2f_AWVALID              : out   std_logic;                                        -- awvalid
			h2f_AWREADY              : in    std_logic                     := 'X';             -- awready
			h2f_WID                  : out   std_logic_vector(11 downto 0);                    -- wid
			h2f_WDATA                : out   std_logic_vector(31 downto 0);                    -- wdata
			h2f_WSTRB                : out   std_logic_vector(3 downto 0);                     -- wstrb
			h2f_WLAST                : out   std_logic;                                        -- wlast
			h2f_WVALID               : out   std_logic;                                        -- wvalid
			h2f_WREADY               : in    std_logic                     := 'X';             -- wready
			h2f_BID                  : in    std_logic_vector(11 downto 0) := (others => 'X'); -- bid
			h2f_BRESP                : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- bresp
			h2f_BVALID               : in    std_logic                     := 'X';             -- bvalid
			h2f_BREADY               : out   std_logic;                                        -- bready
			h2f_ARID                 : out   std_logic_vector(11 downto 0);                    -- arid
			h2f_ARADDR               : out   std_logic_vector(29 downto 0);                    -- araddr
			h2f_ARLEN                : out   std_logic_vector(3 downto 0);                     -- arlen
			h2f_ARSIZE               : out   std_logic_vector(2 downto 0);                     -- arsize
			h2f_ARBURST              : out   std_logic_vector(1 downto 0);                     -- arburst
			h2f_ARLOCK               : out   std_logic_vector(1 downto 0);                     -- arlock
			h2f_ARCACHE              : out   std_logic_vector(3 downto 0);                     -- arcache
			h2f_ARPROT               : out   std_logic_vector(2 downto 0);                     -- arprot
			h2f_ARVALID              : out   std_logic;                                        -- arvalid
			h2f_ARREADY              : in    std_logic                     := 'X';             -- arready
			h2f_RID                  : in    std_logic_vector(11 downto 0) := (others => 'X'); -- rid
			h2f_RDATA                : in    std_logic_vector(31 downto 0) := (others => 'X'); -- rdata
			h2f_RRESP                : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- rresp
			h2f_RLAST                : in    std_logic                     := 'X';             -- rlast
			h2f_RVALID               : in    std_logic                     := 'X';             -- rvalid
			h2f_RREADY               : out   std_logic;                                        -- rready
			f2h_axi_clk              : in    std_logic                     := 'X';             -- clk
			f2h_AWID                 : in    std_logic_vector(7 downto 0)  := (others => 'X'); -- awid
			f2h_AWADDR               : in    std_logic_vector(31 downto 0) := (others => 'X'); -- awaddr
			f2h_AWLEN                : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- awlen
			f2h_AWSIZE               : in    std_logic_vector(2 downto 0)  := (others => 'X'); -- awsize
			f2h_AWBURST              : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- awburst
			f2h_AWLOCK               : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- awlock
			f2h_AWCACHE              : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- awcache
			f2h_AWPROT               : in    std_logic_vector(2 downto 0)  := (others => 'X'); -- awprot
			f2h_AWVALID              : in    std_logic                     := 'X';             -- awvalid
			f2h_AWREADY              : out   std_logic;                                        -- awready
			f2h_AWUSER               : in    std_logic_vector(4 downto 0)  := (others => 'X'); -- awuser
			f2h_WID                  : in    std_logic_vector(7 downto 0)  := (others => 'X'); -- wid
			f2h_WDATA                : in    std_logic_vector(31 downto 0) := (others => 'X'); -- wdata
			f2h_WSTRB                : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- wstrb
			f2h_WLAST                : in    std_logic                     := 'X';             -- wlast
			f2h_WVALID               : in    std_logic                     := 'X';             -- wvalid
			f2h_WREADY               : out   std_logic;                                        -- wready
			f2h_BID                  : out   std_logic_vector(7 downto 0);                     -- bid
			f2h_BRESP                : out   std_logic_vector(1 downto 0);                     -- bresp
			f2h_BVALID               : out   std_logic;                                        -- bvalid
			f2h_BREADY               : in    std_logic                     := 'X';             -- bready
			f2h_ARID                 : in    std_logic_vector(7 downto 0)  := (others => 'X'); -- arid
			f2h_ARADDR               : in    std_logic_vector(31 downto 0) := (others => 'X'); -- araddr
			f2h_ARLEN                : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- arlen
			f2h_ARSIZE               : in    std_logic_vector(2 downto 0)  := (others => 'X'); -- arsize
			f2h_ARBURST              : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- arburst
			f2h_ARLOCK               : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- arlock
			f2h_ARCACHE              : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- arcache
			f2h_ARPROT               : in    std_logic_vector(2 downto 0)  := (others => 'X'); -- arprot
			f2h_ARVALID              : in    std_logic                     := 'X';             -- arvalid
			f2h_ARREADY              : out   std_logic;                                        -- arready
			f2h_ARUSER               : in    std_logic_vector(4 downto 0)  := (others => 'X'); -- aruser
			f2h_RID                  : out   std_logic_vector(7 downto 0);                     -- rid
			f2h_RDATA                : out   std_logic_vector(31 downto 0);                    -- rdata
			f2h_RRESP                : out   std_logic_vector(1 downto 0);                     -- rresp
			f2h_RLAST                : out   std_logic;                                        -- rlast
			f2h_RVALID               : out   std_logic;                                        -- rvalid
			f2h_RREADY               : in    std_logic                     := 'X';             -- rready
			h2f_lw_axi_clk           : in    std_logic                     := 'X';             -- clk
			h2f_lw_AWID              : out   std_logic_vector(11 downto 0);                    -- awid
			h2f_lw_AWADDR            : out   std_logic_vector(20 downto 0);                    -- awaddr
			h2f_lw_AWLEN             : out   std_logic_vector(3 downto 0);                     -- awlen
			h2f_lw_AWSIZE            : out   std_logic_vector(2 downto 0);                     -- awsize
			h2f_lw_AWBURST           : out   std_logic_vector(1 downto 0);                     -- awburst
			h2f_lw_AWLOCK            : out   std_logic_vector(1 downto 0);                     -- awlock
			h2f_lw_AWCACHE           : out   std_logic_vector(3 downto 0);                     -- awcache
			h2f_lw_AWPROT            : out   std_logic_vector(2 downto 0);                     -- awprot
			h2f_lw_AWVALID           : out   std_logic;                                        -- awvalid
			h2f_lw_AWREADY           : in    std_logic                     := 'X';             -- awready
			h2f_lw_WID               : out   std_logic_vector(11 downto 0);                    -- wid
			h2f_lw_WDATA             : out   std_logic_vector(31 downto 0);                    -- wdata
			h2f_lw_WSTRB             : out   std_logic_vector(3 downto 0);                     -- wstrb
			h2f_lw_WLAST             : out   std_logic;                                        -- wlast
			h2f_lw_WVALID            : out   std_logic;                                        -- wvalid
			h2f_lw_WREADY            : in    std_logic                     := 'X';             -- wready
			h2f_lw_BID               : in    std_logic_vector(11 downto 0) := (others => 'X'); -- bid
			h2f_lw_BRESP             : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- bresp
			h2f_lw_BVALID            : in    std_logic                     := 'X';             -- bvalid
			h2f_lw_BREADY            : out   std_logic;                                        -- bready
			h2f_lw_ARID              : out   std_logic_vector(11 downto 0);                    -- arid
			h2f_lw_ARADDR            : out   std_logic_vector(20 downto 0);                    -- araddr
			h2f_lw_ARLEN             : out   std_logic_vector(3 downto 0);                     -- arlen
			h2f_lw_ARSIZE            : out   std_logic_vector(2 downto 0);                     -- arsize
			h2f_lw_ARBURST           : out   std_logic_vector(1 downto 0);                     -- arburst
			h2f_lw_ARLOCK            : out   std_logic_vector(1 downto 0);                     -- arlock
			h2f_lw_ARCACHE           : out   std_logic_vector(3 downto 0);                     -- arcache
			h2f_lw_ARPROT            : out   std_logic_vector(2 downto 0);                     -- arprot
			h2f_lw_ARVALID           : out   std_logic;                                        -- arvalid
			h2f_lw_ARREADY           : in    std_logic                     := 'X';             -- arready
			h2f_lw_RID               : in    std_logic_vector(11 downto 0) := (others => 'X'); -- rid
			h2f_lw_RDATA             : in    std_logic_vector(31 downto 0) := (others => 'X'); -- rdata
			h2f_lw_RRESP             : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- rresp
			h2f_lw_RLAST             : in    std_logic                     := 'X';             -- rlast
			h2f_lw_RVALID            : in    std_logic                     := 'X';             -- rvalid
			h2f_lw_RREADY            : out   std_logic;                                        -- rready
			f2h_irq_p0               : in    std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			f2h_irq_p1               : in    std_logic_vector(31 downto 0) := (others => 'X')  -- irq
		);
	end component standalone_hps_hps_0;

	component standalone_hps_leds_o is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(3 downto 0)                      -- export
		);
	end component standalone_hps_leds_o;

	component standalone_hps_mm_interconnect_0 is
		port (
			axi_bridge_0_s0_awid                               : out std_logic_vector(11 downto 0);                    -- awid
			axi_bridge_0_s0_awaddr                             : out std_logic_vector(29 downto 0);                    -- awaddr
			axi_bridge_0_s0_awlen                              : out std_logic_vector(7 downto 0);                     -- awlen
			axi_bridge_0_s0_awsize                             : out std_logic_vector(2 downto 0);                     -- awsize
			axi_bridge_0_s0_awburst                            : out std_logic_vector(1 downto 0);                     -- awburst
			axi_bridge_0_s0_awlock                             : out std_logic_vector(0 downto 0);                     -- awlock
			axi_bridge_0_s0_awcache                            : out std_logic_vector(3 downto 0);                     -- awcache
			axi_bridge_0_s0_awprot                             : out std_logic_vector(2 downto 0);                     -- awprot
			axi_bridge_0_s0_awqos                              : out std_logic_vector(3 downto 0);                     -- awqos
			axi_bridge_0_s0_awvalid                            : out std_logic;                                        -- awvalid
			axi_bridge_0_s0_awready                            : in  std_logic                     := 'X';             -- awready
			axi_bridge_0_s0_wdata                              : out std_logic_vector(31 downto 0);                    -- wdata
			axi_bridge_0_s0_wstrb                              : out std_logic_vector(3 downto 0);                     -- wstrb
			axi_bridge_0_s0_wlast                              : out std_logic;                                        -- wlast
			axi_bridge_0_s0_wvalid                             : out std_logic;                                        -- wvalid
			axi_bridge_0_s0_wready                             : in  std_logic                     := 'X';             -- wready
			axi_bridge_0_s0_bid                                : in  std_logic_vector(11 downto 0) := (others => 'X'); -- bid
			axi_bridge_0_s0_bresp                              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- bresp
			axi_bridge_0_s0_bvalid                             : in  std_logic                     := 'X';             -- bvalid
			axi_bridge_0_s0_bready                             : out std_logic;                                        -- bready
			axi_bridge_0_s0_arid                               : out std_logic_vector(11 downto 0);                    -- arid
			axi_bridge_0_s0_araddr                             : out std_logic_vector(29 downto 0);                    -- araddr
			axi_bridge_0_s0_arlen                              : out std_logic_vector(7 downto 0);                     -- arlen
			axi_bridge_0_s0_arsize                             : out std_logic_vector(2 downto 0);                     -- arsize
			axi_bridge_0_s0_arburst                            : out std_logic_vector(1 downto 0);                     -- arburst
			axi_bridge_0_s0_arlock                             : out std_logic_vector(0 downto 0);                     -- arlock
			axi_bridge_0_s0_arcache                            : out std_logic_vector(3 downto 0);                     -- arcache
			axi_bridge_0_s0_arprot                             : out std_logic_vector(2 downto 0);                     -- arprot
			axi_bridge_0_s0_arqos                              : out std_logic_vector(3 downto 0);                     -- arqos
			axi_bridge_0_s0_arvalid                            : out std_logic;                                        -- arvalid
			axi_bridge_0_s0_arready                            : in  std_logic                     := 'X';             -- arready
			axi_bridge_0_s0_rid                                : in  std_logic_vector(11 downto 0) := (others => 'X'); -- rid
			axi_bridge_0_s0_rdata                              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- rdata
			axi_bridge_0_s0_rresp                              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- rresp
			axi_bridge_0_s0_rlast                              : in  std_logic                     := 'X';             -- rlast
			axi_bridge_0_s0_rvalid                             : in  std_logic                     := 'X';             -- rvalid
			axi_bridge_0_s0_rready                             : out std_logic;                                        -- rready
			hps_0_h2f_axi_master_awid                          : in  std_logic_vector(11 downto 0) := (others => 'X'); -- awid
			hps_0_h2f_axi_master_awaddr                        : in  std_logic_vector(29 downto 0) := (others => 'X'); -- awaddr
			hps_0_h2f_axi_master_awlen                         : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- awlen
			hps_0_h2f_axi_master_awsize                        : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- awsize
			hps_0_h2f_axi_master_awburst                       : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- awburst
			hps_0_h2f_axi_master_awlock                        : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- awlock
			hps_0_h2f_axi_master_awcache                       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- awcache
			hps_0_h2f_axi_master_awprot                        : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- awprot
			hps_0_h2f_axi_master_awvalid                       : in  std_logic                     := 'X';             -- awvalid
			hps_0_h2f_axi_master_awready                       : out std_logic;                                        -- awready
			hps_0_h2f_axi_master_wid                           : in  std_logic_vector(11 downto 0) := (others => 'X'); -- wid
			hps_0_h2f_axi_master_wdata                         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- wdata
			hps_0_h2f_axi_master_wstrb                         : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- wstrb
			hps_0_h2f_axi_master_wlast                         : in  std_logic                     := 'X';             -- wlast
			hps_0_h2f_axi_master_wvalid                        : in  std_logic                     := 'X';             -- wvalid
			hps_0_h2f_axi_master_wready                        : out std_logic;                                        -- wready
			hps_0_h2f_axi_master_bid                           : out std_logic_vector(11 downto 0);                    -- bid
			hps_0_h2f_axi_master_bresp                         : out std_logic_vector(1 downto 0);                     -- bresp
			hps_0_h2f_axi_master_bvalid                        : out std_logic;                                        -- bvalid
			hps_0_h2f_axi_master_bready                        : in  std_logic                     := 'X';             -- bready
			hps_0_h2f_axi_master_arid                          : in  std_logic_vector(11 downto 0) := (others => 'X'); -- arid
			hps_0_h2f_axi_master_araddr                        : in  std_logic_vector(29 downto 0) := (others => 'X'); -- araddr
			hps_0_h2f_axi_master_arlen                         : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- arlen
			hps_0_h2f_axi_master_arsize                        : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- arsize
			hps_0_h2f_axi_master_arburst                       : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- arburst
			hps_0_h2f_axi_master_arlock                        : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- arlock
			hps_0_h2f_axi_master_arcache                       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- arcache
			hps_0_h2f_axi_master_arprot                        : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- arprot
			hps_0_h2f_axi_master_arvalid                       : in  std_logic                     := 'X';             -- arvalid
			hps_0_h2f_axi_master_arready                       : out std_logic;                                        -- arready
			hps_0_h2f_axi_master_rid                           : out std_logic_vector(11 downto 0);                    -- rid
			hps_0_h2f_axi_master_rdata                         : out std_logic_vector(31 downto 0);                    -- rdata
			hps_0_h2f_axi_master_rresp                         : out std_logic_vector(1 downto 0);                     -- rresp
			hps_0_h2f_axi_master_rlast                         : out std_logic;                                        -- rlast
			hps_0_h2f_axi_master_rvalid                        : out std_logic;                                        -- rvalid
			hps_0_h2f_axi_master_rready                        : in  std_logic                     := 'X';             -- rready
			clk_0_clk_clk                                      : in  std_logic                     := 'X';             -- clk
			axi_bridge_0_clk_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X'              -- reset
		);
	end component standalone_hps_mm_interconnect_0;

	component standalone_hps_mm_interconnect_1 is
		port (
			hps_0_h2f_lw_axi_master_awid                                        : in  std_logic_vector(11 downto 0) := (others => 'X'); -- awid
			hps_0_h2f_lw_axi_master_awaddr                                      : in  std_logic_vector(20 downto 0) := (others => 'X'); -- awaddr
			hps_0_h2f_lw_axi_master_awlen                                       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- awlen
			hps_0_h2f_lw_axi_master_awsize                                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- awsize
			hps_0_h2f_lw_axi_master_awburst                                     : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- awburst
			hps_0_h2f_lw_axi_master_awlock                                      : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- awlock
			hps_0_h2f_lw_axi_master_awcache                                     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- awcache
			hps_0_h2f_lw_axi_master_awprot                                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- awprot
			hps_0_h2f_lw_axi_master_awvalid                                     : in  std_logic                     := 'X';             -- awvalid
			hps_0_h2f_lw_axi_master_awready                                     : out std_logic;                                        -- awready
			hps_0_h2f_lw_axi_master_wid                                         : in  std_logic_vector(11 downto 0) := (others => 'X'); -- wid
			hps_0_h2f_lw_axi_master_wdata                                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- wdata
			hps_0_h2f_lw_axi_master_wstrb                                       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- wstrb
			hps_0_h2f_lw_axi_master_wlast                                       : in  std_logic                     := 'X';             -- wlast
			hps_0_h2f_lw_axi_master_wvalid                                      : in  std_logic                     := 'X';             -- wvalid
			hps_0_h2f_lw_axi_master_wready                                      : out std_logic;                                        -- wready
			hps_0_h2f_lw_axi_master_bid                                         : out std_logic_vector(11 downto 0);                    -- bid
			hps_0_h2f_lw_axi_master_bresp                                       : out std_logic_vector(1 downto 0);                     -- bresp
			hps_0_h2f_lw_axi_master_bvalid                                      : out std_logic;                                        -- bvalid
			hps_0_h2f_lw_axi_master_bready                                      : in  std_logic                     := 'X';             -- bready
			hps_0_h2f_lw_axi_master_arid                                        : in  std_logic_vector(11 downto 0) := (others => 'X'); -- arid
			hps_0_h2f_lw_axi_master_araddr                                      : in  std_logic_vector(20 downto 0) := (others => 'X'); -- araddr
			hps_0_h2f_lw_axi_master_arlen                                       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- arlen
			hps_0_h2f_lw_axi_master_arsize                                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- arsize
			hps_0_h2f_lw_axi_master_arburst                                     : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- arburst
			hps_0_h2f_lw_axi_master_arlock                                      : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- arlock
			hps_0_h2f_lw_axi_master_arcache                                     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- arcache
			hps_0_h2f_lw_axi_master_arprot                                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- arprot
			hps_0_h2f_lw_axi_master_arvalid                                     : in  std_logic                     := 'X';             -- arvalid
			hps_0_h2f_lw_axi_master_arready                                     : out std_logic;                                        -- arready
			hps_0_h2f_lw_axi_master_rid                                         : out std_logic_vector(11 downto 0);                    -- rid
			hps_0_h2f_lw_axi_master_rdata                                       : out std_logic_vector(31 downto 0);                    -- rdata
			hps_0_h2f_lw_axi_master_rresp                                       : out std_logic_vector(1 downto 0);                     -- rresp
			hps_0_h2f_lw_axi_master_rlast                                       : out std_logic;                                        -- rlast
			hps_0_h2f_lw_axi_master_rvalid                                      : out std_logic;                                        -- rvalid
			hps_0_h2f_lw_axi_master_rready                                      : in  std_logic                     := 'X';             -- rready
			clk_0_clk_clk                                                       : in  std_logic                     := 'X';             -- clk
			hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			leds_o_reset_reset_bridge_in_reset_reset                            : in  std_logic                     := 'X';             -- reset
			buttons_i_s1_address                                                : out std_logic_vector(1 downto 0);                     -- address
			buttons_i_s1_readdata                                               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			dipsw_i_s1_address                                                  : out std_logic_vector(1 downto 0);                     -- address
			dipsw_i_s1_readdata                                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			leds_o_s1_address                                                   : out std_logic_vector(1 downto 0);                     -- address
			leds_o_s1_write                                                     : out std_logic;                                        -- write
			leds_o_s1_readdata                                                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			leds_o_s1_writedata                                                 : out std_logic_vector(31 downto 0);                    -- writedata
			leds_o_s1_chipselect                                                : out std_logic                                         -- chipselect
		);
	end component standalone_hps_mm_interconnect_1;

	component standalone_hps_irq_mapper is
		port (
			clk        : in  std_logic                     := 'X'; -- clk
			reset      : in  std_logic                     := 'X'; -- reset
			sender_irq : out std_logic_vector(31 downto 0)         -- irq
		);
	end component standalone_hps_irq_mapper;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	signal hps_0_h2f_reset_reset                       : std_logic;                     -- hps_0:h2f_rst_n -> [h2f_reset_reset_n, h2f_reset_reset_n:in]
	signal hps_0_h2f_axi_master_awburst                : std_logic_vector(1 downto 0);  -- hps_0:h2f_AWBURST -> mm_interconnect_0:hps_0_h2f_axi_master_awburst
	signal hps_0_h2f_axi_master_arlen                  : std_logic_vector(3 downto 0);  -- hps_0:h2f_ARLEN -> mm_interconnect_0:hps_0_h2f_axi_master_arlen
	signal hps_0_h2f_axi_master_wstrb                  : std_logic_vector(3 downto 0);  -- hps_0:h2f_WSTRB -> mm_interconnect_0:hps_0_h2f_axi_master_wstrb
	signal hps_0_h2f_axi_master_wready                 : std_logic;                     -- mm_interconnect_0:hps_0_h2f_axi_master_wready -> hps_0:h2f_WREADY
	signal hps_0_h2f_axi_master_rid                    : std_logic_vector(11 downto 0); -- mm_interconnect_0:hps_0_h2f_axi_master_rid -> hps_0:h2f_RID
	signal hps_0_h2f_axi_master_rready                 : std_logic;                     -- hps_0:h2f_RREADY -> mm_interconnect_0:hps_0_h2f_axi_master_rready
	signal hps_0_h2f_axi_master_awlen                  : std_logic_vector(3 downto 0);  -- hps_0:h2f_AWLEN -> mm_interconnect_0:hps_0_h2f_axi_master_awlen
	signal hps_0_h2f_axi_master_wid                    : std_logic_vector(11 downto 0); -- hps_0:h2f_WID -> mm_interconnect_0:hps_0_h2f_axi_master_wid
	signal hps_0_h2f_axi_master_arcache                : std_logic_vector(3 downto 0);  -- hps_0:h2f_ARCACHE -> mm_interconnect_0:hps_0_h2f_axi_master_arcache
	signal hps_0_h2f_axi_master_wvalid                 : std_logic;                     -- hps_0:h2f_WVALID -> mm_interconnect_0:hps_0_h2f_axi_master_wvalid
	signal hps_0_h2f_axi_master_araddr                 : std_logic_vector(29 downto 0); -- hps_0:h2f_ARADDR -> mm_interconnect_0:hps_0_h2f_axi_master_araddr
	signal hps_0_h2f_axi_master_arprot                 : std_logic_vector(2 downto 0);  -- hps_0:h2f_ARPROT -> mm_interconnect_0:hps_0_h2f_axi_master_arprot
	signal hps_0_h2f_axi_master_awprot                 : std_logic_vector(2 downto 0);  -- hps_0:h2f_AWPROT -> mm_interconnect_0:hps_0_h2f_axi_master_awprot
	signal hps_0_h2f_axi_master_wdata                  : std_logic_vector(31 downto 0); -- hps_0:h2f_WDATA -> mm_interconnect_0:hps_0_h2f_axi_master_wdata
	signal hps_0_h2f_axi_master_arvalid                : std_logic;                     -- hps_0:h2f_ARVALID -> mm_interconnect_0:hps_0_h2f_axi_master_arvalid
	signal hps_0_h2f_axi_master_awcache                : std_logic_vector(3 downto 0);  -- hps_0:h2f_AWCACHE -> mm_interconnect_0:hps_0_h2f_axi_master_awcache
	signal hps_0_h2f_axi_master_arid                   : std_logic_vector(11 downto 0); -- hps_0:h2f_ARID -> mm_interconnect_0:hps_0_h2f_axi_master_arid
	signal hps_0_h2f_axi_master_arlock                 : std_logic_vector(1 downto 0);  -- hps_0:h2f_ARLOCK -> mm_interconnect_0:hps_0_h2f_axi_master_arlock
	signal hps_0_h2f_axi_master_awlock                 : std_logic_vector(1 downto 0);  -- hps_0:h2f_AWLOCK -> mm_interconnect_0:hps_0_h2f_axi_master_awlock
	signal hps_0_h2f_axi_master_awaddr                 : std_logic_vector(29 downto 0); -- hps_0:h2f_AWADDR -> mm_interconnect_0:hps_0_h2f_axi_master_awaddr
	signal hps_0_h2f_axi_master_bresp                  : std_logic_vector(1 downto 0);  -- mm_interconnect_0:hps_0_h2f_axi_master_bresp -> hps_0:h2f_BRESP
	signal hps_0_h2f_axi_master_arready                : std_logic;                     -- mm_interconnect_0:hps_0_h2f_axi_master_arready -> hps_0:h2f_ARREADY
	signal hps_0_h2f_axi_master_rdata                  : std_logic_vector(31 downto 0); -- mm_interconnect_0:hps_0_h2f_axi_master_rdata -> hps_0:h2f_RDATA
	signal hps_0_h2f_axi_master_awready                : std_logic;                     -- mm_interconnect_0:hps_0_h2f_axi_master_awready -> hps_0:h2f_AWREADY
	signal hps_0_h2f_axi_master_arburst                : std_logic_vector(1 downto 0);  -- hps_0:h2f_ARBURST -> mm_interconnect_0:hps_0_h2f_axi_master_arburst
	signal hps_0_h2f_axi_master_arsize                 : std_logic_vector(2 downto 0);  -- hps_0:h2f_ARSIZE -> mm_interconnect_0:hps_0_h2f_axi_master_arsize
	signal hps_0_h2f_axi_master_bready                 : std_logic;                     -- hps_0:h2f_BREADY -> mm_interconnect_0:hps_0_h2f_axi_master_bready
	signal hps_0_h2f_axi_master_rlast                  : std_logic;                     -- mm_interconnect_0:hps_0_h2f_axi_master_rlast -> hps_0:h2f_RLAST
	signal hps_0_h2f_axi_master_wlast                  : std_logic;                     -- hps_0:h2f_WLAST -> mm_interconnect_0:hps_0_h2f_axi_master_wlast
	signal hps_0_h2f_axi_master_rresp                  : std_logic_vector(1 downto 0);  -- mm_interconnect_0:hps_0_h2f_axi_master_rresp -> hps_0:h2f_RRESP
	signal hps_0_h2f_axi_master_awid                   : std_logic_vector(11 downto 0); -- hps_0:h2f_AWID -> mm_interconnect_0:hps_0_h2f_axi_master_awid
	signal hps_0_h2f_axi_master_bid                    : std_logic_vector(11 downto 0); -- mm_interconnect_0:hps_0_h2f_axi_master_bid -> hps_0:h2f_BID
	signal hps_0_h2f_axi_master_bvalid                 : std_logic;                     -- mm_interconnect_0:hps_0_h2f_axi_master_bvalid -> hps_0:h2f_BVALID
	signal hps_0_h2f_axi_master_awsize                 : std_logic_vector(2 downto 0);  -- hps_0:h2f_AWSIZE -> mm_interconnect_0:hps_0_h2f_axi_master_awsize
	signal hps_0_h2f_axi_master_awvalid                : std_logic;                     -- hps_0:h2f_AWVALID -> mm_interconnect_0:hps_0_h2f_axi_master_awvalid
	signal hps_0_h2f_axi_master_rvalid                 : std_logic;                     -- mm_interconnect_0:hps_0_h2f_axi_master_rvalid -> hps_0:h2f_RVALID
	signal mm_interconnect_0_axi_bridge_0_s0_awburst   : std_logic_vector(1 downto 0);  -- mm_interconnect_0:axi_bridge_0_s0_awburst -> axi_bridge_0:s0_awburst
	signal mm_interconnect_0_axi_bridge_0_s0_arlen     : std_logic_vector(7 downto 0);  -- mm_interconnect_0:axi_bridge_0_s0_arlen -> axi_bridge_0:s0_arlen
	signal mm_interconnect_0_axi_bridge_0_s0_arqos     : std_logic_vector(3 downto 0);  -- mm_interconnect_0:axi_bridge_0_s0_arqos -> axi_bridge_0:s0_arqos
	signal mm_interconnect_0_axi_bridge_0_s0_wstrb     : std_logic_vector(3 downto 0);  -- mm_interconnect_0:axi_bridge_0_s0_wstrb -> axi_bridge_0:s0_wstrb
	signal mm_interconnect_0_axi_bridge_0_s0_wready    : std_logic;                     -- axi_bridge_0:s0_wready -> mm_interconnect_0:axi_bridge_0_s0_wready
	signal mm_interconnect_0_axi_bridge_0_s0_rid       : std_logic_vector(11 downto 0); -- axi_bridge_0:s0_rid -> mm_interconnect_0:axi_bridge_0_s0_rid
	signal mm_interconnect_0_axi_bridge_0_s0_rready    : std_logic;                     -- mm_interconnect_0:axi_bridge_0_s0_rready -> axi_bridge_0:s0_rready
	signal mm_interconnect_0_axi_bridge_0_s0_awlen     : std_logic_vector(7 downto 0);  -- mm_interconnect_0:axi_bridge_0_s0_awlen -> axi_bridge_0:s0_awlen
	signal mm_interconnect_0_axi_bridge_0_s0_awqos     : std_logic_vector(3 downto 0);  -- mm_interconnect_0:axi_bridge_0_s0_awqos -> axi_bridge_0:s0_awqos
	signal mm_interconnect_0_axi_bridge_0_s0_arcache   : std_logic_vector(3 downto 0);  -- mm_interconnect_0:axi_bridge_0_s0_arcache -> axi_bridge_0:s0_arcache
	signal mm_interconnect_0_axi_bridge_0_s0_wvalid    : std_logic;                     -- mm_interconnect_0:axi_bridge_0_s0_wvalid -> axi_bridge_0:s0_wvalid
	signal mm_interconnect_0_axi_bridge_0_s0_araddr    : std_logic_vector(29 downto 0); -- mm_interconnect_0:axi_bridge_0_s0_araddr -> axi_bridge_0:s0_araddr
	signal mm_interconnect_0_axi_bridge_0_s0_arprot    : std_logic_vector(2 downto 0);  -- mm_interconnect_0:axi_bridge_0_s0_arprot -> axi_bridge_0:s0_arprot
	signal mm_interconnect_0_axi_bridge_0_s0_awprot    : std_logic_vector(2 downto 0);  -- mm_interconnect_0:axi_bridge_0_s0_awprot -> axi_bridge_0:s0_awprot
	signal mm_interconnect_0_axi_bridge_0_s0_wdata     : std_logic_vector(31 downto 0); -- mm_interconnect_0:axi_bridge_0_s0_wdata -> axi_bridge_0:s0_wdata
	signal mm_interconnect_0_axi_bridge_0_s0_arvalid   : std_logic;                     -- mm_interconnect_0:axi_bridge_0_s0_arvalid -> axi_bridge_0:s0_arvalid
	signal mm_interconnect_0_axi_bridge_0_s0_awcache   : std_logic_vector(3 downto 0);  -- mm_interconnect_0:axi_bridge_0_s0_awcache -> axi_bridge_0:s0_awcache
	signal mm_interconnect_0_axi_bridge_0_s0_arid      : std_logic_vector(11 downto 0); -- mm_interconnect_0:axi_bridge_0_s0_arid -> axi_bridge_0:s0_arid
	signal mm_interconnect_0_axi_bridge_0_s0_arlock    : std_logic_vector(0 downto 0);  -- mm_interconnect_0:axi_bridge_0_s0_arlock -> axi_bridge_0:s0_arlock
	signal mm_interconnect_0_axi_bridge_0_s0_awlock    : std_logic_vector(0 downto 0);  -- mm_interconnect_0:axi_bridge_0_s0_awlock -> axi_bridge_0:s0_awlock
	signal mm_interconnect_0_axi_bridge_0_s0_awaddr    : std_logic_vector(29 downto 0); -- mm_interconnect_0:axi_bridge_0_s0_awaddr -> axi_bridge_0:s0_awaddr
	signal mm_interconnect_0_axi_bridge_0_s0_bresp     : std_logic_vector(1 downto 0);  -- axi_bridge_0:s0_bresp -> mm_interconnect_0:axi_bridge_0_s0_bresp
	signal mm_interconnect_0_axi_bridge_0_s0_arready   : std_logic;                     -- axi_bridge_0:s0_arready -> mm_interconnect_0:axi_bridge_0_s0_arready
	signal mm_interconnect_0_axi_bridge_0_s0_rdata     : std_logic_vector(31 downto 0); -- axi_bridge_0:s0_rdata -> mm_interconnect_0:axi_bridge_0_s0_rdata
	signal mm_interconnect_0_axi_bridge_0_s0_awready   : std_logic;                     -- axi_bridge_0:s0_awready -> mm_interconnect_0:axi_bridge_0_s0_awready
	signal mm_interconnect_0_axi_bridge_0_s0_arburst   : std_logic_vector(1 downto 0);  -- mm_interconnect_0:axi_bridge_0_s0_arburst -> axi_bridge_0:s0_arburst
	signal mm_interconnect_0_axi_bridge_0_s0_arsize    : std_logic_vector(2 downto 0);  -- mm_interconnect_0:axi_bridge_0_s0_arsize -> axi_bridge_0:s0_arsize
	signal mm_interconnect_0_axi_bridge_0_s0_bready    : std_logic;                     -- mm_interconnect_0:axi_bridge_0_s0_bready -> axi_bridge_0:s0_bready
	signal mm_interconnect_0_axi_bridge_0_s0_rlast     : std_logic;                     -- axi_bridge_0:s0_rlast -> mm_interconnect_0:axi_bridge_0_s0_rlast
	signal mm_interconnect_0_axi_bridge_0_s0_wlast     : std_logic;                     -- mm_interconnect_0:axi_bridge_0_s0_wlast -> axi_bridge_0:s0_wlast
	signal mm_interconnect_0_axi_bridge_0_s0_rresp     : std_logic_vector(1 downto 0);  -- axi_bridge_0:s0_rresp -> mm_interconnect_0:axi_bridge_0_s0_rresp
	signal mm_interconnect_0_axi_bridge_0_s0_awid      : std_logic_vector(11 downto 0); -- mm_interconnect_0:axi_bridge_0_s0_awid -> axi_bridge_0:s0_awid
	signal mm_interconnect_0_axi_bridge_0_s0_bid       : std_logic_vector(11 downto 0); -- axi_bridge_0:s0_bid -> mm_interconnect_0:axi_bridge_0_s0_bid
	signal mm_interconnect_0_axi_bridge_0_s0_bvalid    : std_logic;                     -- axi_bridge_0:s0_bvalid -> mm_interconnect_0:axi_bridge_0_s0_bvalid
	signal mm_interconnect_0_axi_bridge_0_s0_awsize    : std_logic_vector(2 downto 0);  -- mm_interconnect_0:axi_bridge_0_s0_awsize -> axi_bridge_0:s0_awsize
	signal mm_interconnect_0_axi_bridge_0_s0_awvalid   : std_logic;                     -- mm_interconnect_0:axi_bridge_0_s0_awvalid -> axi_bridge_0:s0_awvalid
	signal mm_interconnect_0_axi_bridge_0_s0_rvalid    : std_logic;                     -- axi_bridge_0:s0_rvalid -> mm_interconnect_0:axi_bridge_0_s0_rvalid
	signal hps_0_h2f_lw_axi_master_awburst             : std_logic_vector(1 downto 0);  -- hps_0:h2f_lw_AWBURST -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awburst
	signal hps_0_h2f_lw_axi_master_arlen               : std_logic_vector(3 downto 0);  -- hps_0:h2f_lw_ARLEN -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arlen
	signal hps_0_h2f_lw_axi_master_wstrb               : std_logic_vector(3 downto 0);  -- hps_0:h2f_lw_WSTRB -> mm_interconnect_1:hps_0_h2f_lw_axi_master_wstrb
	signal hps_0_h2f_lw_axi_master_wready              : std_logic;                     -- mm_interconnect_1:hps_0_h2f_lw_axi_master_wready -> hps_0:h2f_lw_WREADY
	signal hps_0_h2f_lw_axi_master_rid                 : std_logic_vector(11 downto 0); -- mm_interconnect_1:hps_0_h2f_lw_axi_master_rid -> hps_0:h2f_lw_RID
	signal hps_0_h2f_lw_axi_master_rready              : std_logic;                     -- hps_0:h2f_lw_RREADY -> mm_interconnect_1:hps_0_h2f_lw_axi_master_rready
	signal hps_0_h2f_lw_axi_master_awlen               : std_logic_vector(3 downto 0);  -- hps_0:h2f_lw_AWLEN -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awlen
	signal hps_0_h2f_lw_axi_master_wid                 : std_logic_vector(11 downto 0); -- hps_0:h2f_lw_WID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_wid
	signal hps_0_h2f_lw_axi_master_arcache             : std_logic_vector(3 downto 0);  -- hps_0:h2f_lw_ARCACHE -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arcache
	signal hps_0_h2f_lw_axi_master_wvalid              : std_logic;                     -- hps_0:h2f_lw_WVALID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_wvalid
	signal hps_0_h2f_lw_axi_master_araddr              : std_logic_vector(20 downto 0); -- hps_0:h2f_lw_ARADDR -> mm_interconnect_1:hps_0_h2f_lw_axi_master_araddr
	signal hps_0_h2f_lw_axi_master_arprot              : std_logic_vector(2 downto 0);  -- hps_0:h2f_lw_ARPROT -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arprot
	signal hps_0_h2f_lw_axi_master_awprot              : std_logic_vector(2 downto 0);  -- hps_0:h2f_lw_AWPROT -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awprot
	signal hps_0_h2f_lw_axi_master_wdata               : std_logic_vector(31 downto 0); -- hps_0:h2f_lw_WDATA -> mm_interconnect_1:hps_0_h2f_lw_axi_master_wdata
	signal hps_0_h2f_lw_axi_master_arvalid             : std_logic;                     -- hps_0:h2f_lw_ARVALID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arvalid
	signal hps_0_h2f_lw_axi_master_awcache             : std_logic_vector(3 downto 0);  -- hps_0:h2f_lw_AWCACHE -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awcache
	signal hps_0_h2f_lw_axi_master_arid                : std_logic_vector(11 downto 0); -- hps_0:h2f_lw_ARID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arid
	signal hps_0_h2f_lw_axi_master_arlock              : std_logic_vector(1 downto 0);  -- hps_0:h2f_lw_ARLOCK -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arlock
	signal hps_0_h2f_lw_axi_master_awlock              : std_logic_vector(1 downto 0);  -- hps_0:h2f_lw_AWLOCK -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awlock
	signal hps_0_h2f_lw_axi_master_awaddr              : std_logic_vector(20 downto 0); -- hps_0:h2f_lw_AWADDR -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awaddr
	signal hps_0_h2f_lw_axi_master_bresp               : std_logic_vector(1 downto 0);  -- mm_interconnect_1:hps_0_h2f_lw_axi_master_bresp -> hps_0:h2f_lw_BRESP
	signal hps_0_h2f_lw_axi_master_arready             : std_logic;                     -- mm_interconnect_1:hps_0_h2f_lw_axi_master_arready -> hps_0:h2f_lw_ARREADY
	signal hps_0_h2f_lw_axi_master_rdata               : std_logic_vector(31 downto 0); -- mm_interconnect_1:hps_0_h2f_lw_axi_master_rdata -> hps_0:h2f_lw_RDATA
	signal hps_0_h2f_lw_axi_master_awready             : std_logic;                     -- mm_interconnect_1:hps_0_h2f_lw_axi_master_awready -> hps_0:h2f_lw_AWREADY
	signal hps_0_h2f_lw_axi_master_arburst             : std_logic_vector(1 downto 0);  -- hps_0:h2f_lw_ARBURST -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arburst
	signal hps_0_h2f_lw_axi_master_arsize              : std_logic_vector(2 downto 0);  -- hps_0:h2f_lw_ARSIZE -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arsize
	signal hps_0_h2f_lw_axi_master_bready              : std_logic;                     -- hps_0:h2f_lw_BREADY -> mm_interconnect_1:hps_0_h2f_lw_axi_master_bready
	signal hps_0_h2f_lw_axi_master_rlast               : std_logic;                     -- mm_interconnect_1:hps_0_h2f_lw_axi_master_rlast -> hps_0:h2f_lw_RLAST
	signal hps_0_h2f_lw_axi_master_wlast               : std_logic;                     -- hps_0:h2f_lw_WLAST -> mm_interconnect_1:hps_0_h2f_lw_axi_master_wlast
	signal hps_0_h2f_lw_axi_master_rresp               : std_logic_vector(1 downto 0);  -- mm_interconnect_1:hps_0_h2f_lw_axi_master_rresp -> hps_0:h2f_lw_RRESP
	signal hps_0_h2f_lw_axi_master_awid                : std_logic_vector(11 downto 0); -- hps_0:h2f_lw_AWID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awid
	signal hps_0_h2f_lw_axi_master_bid                 : std_logic_vector(11 downto 0); -- mm_interconnect_1:hps_0_h2f_lw_axi_master_bid -> hps_0:h2f_lw_BID
	signal hps_0_h2f_lw_axi_master_bvalid              : std_logic;                     -- mm_interconnect_1:hps_0_h2f_lw_axi_master_bvalid -> hps_0:h2f_lw_BVALID
	signal hps_0_h2f_lw_axi_master_awsize              : std_logic_vector(2 downto 0);  -- hps_0:h2f_lw_AWSIZE -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awsize
	signal hps_0_h2f_lw_axi_master_awvalid             : std_logic;                     -- hps_0:h2f_lw_AWVALID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awvalid
	signal hps_0_h2f_lw_axi_master_rvalid              : std_logic;                     -- mm_interconnect_1:hps_0_h2f_lw_axi_master_rvalid -> hps_0:h2f_lw_RVALID
	signal mm_interconnect_1_leds_o_s1_chipselect      : std_logic;                     -- mm_interconnect_1:leds_o_s1_chipselect -> leds_o:chipselect
	signal mm_interconnect_1_leds_o_s1_readdata        : std_logic_vector(31 downto 0); -- leds_o:readdata -> mm_interconnect_1:leds_o_s1_readdata
	signal mm_interconnect_1_leds_o_s1_address         : std_logic_vector(1 downto 0);  -- mm_interconnect_1:leds_o_s1_address -> leds_o:address
	signal mm_interconnect_1_leds_o_s1_write           : std_logic;                     -- mm_interconnect_1:leds_o_s1_write -> mm_interconnect_1_leds_o_s1_write:in
	signal mm_interconnect_1_leds_o_s1_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_1:leds_o_s1_writedata -> leds_o:writedata
	signal mm_interconnect_1_dipsw_i_s1_readdata       : std_logic_vector(31 downto 0); -- dipsw_i:readdata -> mm_interconnect_1:dipsw_i_s1_readdata
	signal mm_interconnect_1_dipsw_i_s1_address        : std_logic_vector(1 downto 0);  -- mm_interconnect_1:dipsw_i_s1_address -> dipsw_i:address
	signal mm_interconnect_1_buttons_i_s1_readdata     : std_logic_vector(31 downto 0); -- buttons_i:readdata -> mm_interconnect_1:buttons_i_s1_readdata
	signal mm_interconnect_1_buttons_i_s1_address      : std_logic_vector(1 downto 0);  -- mm_interconnect_1:buttons_i_s1_address -> buttons_i:address
	signal hps_0_f2h_irq0_irq                          : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> hps_0:f2h_irq_p0
	signal hps_0_f2h_irq1_irq                          : std_logic_vector(31 downto 0); -- irq_mapper_001:sender_irq -> hps_0:f2h_irq_p1
	signal rst_controller_reset_out_reset              : std_logic;                     -- rst_controller:reset_out -> [mm_interconnect_0:axi_bridge_0_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_1:leds_o_reset_reset_bridge_in_reset_reset, rst_controller_reset_out_reset:in]
	signal rst_controller_001_reset_out_reset          : std_logic;                     -- rst_controller_001:reset_out -> mm_interconnect_1:hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset
	signal h2f_reset_reset_n_ports_inv                 : std_logic;                     -- h2f_reset_reset_n:inv -> rst_controller_001:reset_in0
	signal reset_reset_n_ports_inv                     : std_logic;                     -- reset_reset_n:inv -> rst_controller:reset_in0
	signal mm_interconnect_1_leds_o_s1_write_ports_inv : std_logic;                     -- mm_interconnect_1_leds_o_s1_write:inv -> leds_o:write_n
	signal rst_controller_reset_out_reset_ports_inv    : std_logic;                     -- rst_controller_reset_out_reset:inv -> [axi_bridge_0:aresetn, buttons_i:reset_n, dipsw_i:reset_n, leds_o:reset_n]

begin

	axi_bridge_0 : component altera_axi_bridge
		generic map (
			USE_PIPELINE          => 1,
			USE_M0_AWID           => 1,
			USE_M0_AWREGION       => 0,
			USE_M0_AWLEN          => 1,
			USE_M0_AWSIZE         => 1,
			USE_M0_AWBURST        => 1,
			USE_M0_AWLOCK         => 1,
			USE_M0_AWCACHE        => 1,
			USE_M0_AWQOS          => 1,
			USE_S0_AWREGION       => 0,
			USE_S0_AWLOCK         => 1,
			USE_S0_AWCACHE        => 1,
			USE_S0_AWQOS          => 1,
			USE_S0_AWPROT         => 1,
			USE_M0_WSTRB          => 1,
			USE_S0_WLAST          => 1,
			USE_M0_BID            => 1,
			USE_M0_BRESP          => 1,
			USE_S0_BRESP          => 1,
			USE_M0_ARID           => 1,
			USE_M0_ARREGION       => 0,
			USE_M0_ARLEN          => 1,
			USE_M0_ARSIZE         => 1,
			USE_M0_ARBURST        => 1,
			USE_M0_ARLOCK         => 1,
			USE_M0_ARCACHE        => 1,
			USE_M0_ARQOS          => 1,
			USE_S0_ARREGION       => 0,
			USE_S0_ARLOCK         => 1,
			USE_S0_ARCACHE        => 1,
			USE_S0_ARQOS          => 1,
			USE_S0_ARPROT         => 1,
			USE_M0_RID            => 1,
			USE_M0_RRESP          => 1,
			USE_M0_RLAST          => 1,
			USE_S0_RRESP          => 1,
			M0_ID_WIDTH           => 12,
			S0_ID_WIDTH           => 12,
			DATA_WIDTH            => 32,
			WRITE_ADDR_USER_WIDTH => 64,
			READ_ADDR_USER_WIDTH  => 64,
			WRITE_DATA_USER_WIDTH => 64,
			WRITE_RESP_USER_WIDTH => 64,
			READ_DATA_USER_WIDTH  => 64,
			ADDR_WIDTH            => 30,
			USE_S0_AWUSER         => 0,
			USE_S0_ARUSER         => 0,
			USE_S0_WUSER          => 0,
			USE_S0_RUSER          => 0,
			USE_S0_BUSER          => 0,
			USE_M0_AWUSER         => 0,
			USE_M0_ARUSER         => 0,
			USE_M0_WUSER          => 0,
			USE_M0_RUSER          => 0,
			USE_M0_BUSER          => 0,
			AXI_VERSION           => "AXI4",
			BURST_LENGTH_WIDTH    => 8,
			LOCK_WIDTH            => 1
		)
		port map (
			aclk        => clk_clk,                                                            --       clk.clk
			aresetn     => rst_controller_reset_out_reset_ports_inv,                           -- clk_reset.reset_n
			s0_awid     => mm_interconnect_0_axi_bridge_0_s0_awid,                             --        s0.awid
			s0_awaddr   => mm_interconnect_0_axi_bridge_0_s0_awaddr,                           --          .awaddr
			s0_awlen    => mm_interconnect_0_axi_bridge_0_s0_awlen,                            --          .awlen
			s0_awsize   => mm_interconnect_0_axi_bridge_0_s0_awsize,                           --          .awsize
			s0_awburst  => mm_interconnect_0_axi_bridge_0_s0_awburst,                          --          .awburst
			s0_awlock   => mm_interconnect_0_axi_bridge_0_s0_awlock,                           --          .awlock
			s0_awcache  => mm_interconnect_0_axi_bridge_0_s0_awcache,                          --          .awcache
			s0_awprot   => mm_interconnect_0_axi_bridge_0_s0_awprot,                           --          .awprot
			s0_awqos    => mm_interconnect_0_axi_bridge_0_s0_awqos,                            --          .awqos
			s0_awvalid  => mm_interconnect_0_axi_bridge_0_s0_awvalid,                          --          .awvalid
			s0_awready  => mm_interconnect_0_axi_bridge_0_s0_awready,                          --          .awready
			s0_wdata    => mm_interconnect_0_axi_bridge_0_s0_wdata,                            --          .wdata
			s0_wstrb    => mm_interconnect_0_axi_bridge_0_s0_wstrb,                            --          .wstrb
			s0_wlast    => mm_interconnect_0_axi_bridge_0_s0_wlast,                            --          .wlast
			s0_wvalid   => mm_interconnect_0_axi_bridge_0_s0_wvalid,                           --          .wvalid
			s0_wready   => mm_interconnect_0_axi_bridge_0_s0_wready,                           --          .wready
			s0_bid      => mm_interconnect_0_axi_bridge_0_s0_bid,                              --          .bid
			s0_bresp    => mm_interconnect_0_axi_bridge_0_s0_bresp,                            --          .bresp
			s0_bvalid   => mm_interconnect_0_axi_bridge_0_s0_bvalid,                           --          .bvalid
			s0_bready   => mm_interconnect_0_axi_bridge_0_s0_bready,                           --          .bready
			s0_arid     => mm_interconnect_0_axi_bridge_0_s0_arid,                             --          .arid
			s0_araddr   => mm_interconnect_0_axi_bridge_0_s0_araddr,                           --          .araddr
			s0_arlen    => mm_interconnect_0_axi_bridge_0_s0_arlen,                            --          .arlen
			s0_arsize   => mm_interconnect_0_axi_bridge_0_s0_arsize,                           --          .arsize
			s0_arburst  => mm_interconnect_0_axi_bridge_0_s0_arburst,                          --          .arburst
			s0_arlock   => mm_interconnect_0_axi_bridge_0_s0_arlock,                           --          .arlock
			s0_arcache  => mm_interconnect_0_axi_bridge_0_s0_arcache,                          --          .arcache
			s0_arprot   => mm_interconnect_0_axi_bridge_0_s0_arprot,                           --          .arprot
			s0_arqos    => mm_interconnect_0_axi_bridge_0_s0_arqos,                            --          .arqos
			s0_arvalid  => mm_interconnect_0_axi_bridge_0_s0_arvalid,                          --          .arvalid
			s0_arready  => mm_interconnect_0_axi_bridge_0_s0_arready,                          --          .arready
			s0_rid      => mm_interconnect_0_axi_bridge_0_s0_rid,                              --          .rid
			s0_rdata    => mm_interconnect_0_axi_bridge_0_s0_rdata,                            --          .rdata
			s0_rresp    => mm_interconnect_0_axi_bridge_0_s0_rresp,                            --          .rresp
			s0_rlast    => mm_interconnect_0_axi_bridge_0_s0_rlast,                            --          .rlast
			s0_rvalid   => mm_interconnect_0_axi_bridge_0_s0_rvalid,                           --          .rvalid
			s0_rready   => mm_interconnect_0_axi_bridge_0_s0_rready,                           --          .rready
			m0_awid     => h2f_bus_awid,                                                       --        m0.awid
			m0_awaddr   => h2f_bus_awaddr,                                                     --          .awaddr
			m0_awlen    => h2f_bus_awlen,                                                      --          .awlen
			m0_awsize   => h2f_bus_awsize,                                                     --          .awsize
			m0_awburst  => h2f_bus_awburst,                                                    --          .awburst
			m0_awlock   => h2f_bus_awlock,                                                     --          .awlock
			m0_awcache  => h2f_bus_awcache,                                                    --          .awcache
			m0_awprot   => h2f_bus_awprot,                                                     --          .awprot
			m0_awqos    => h2f_bus_awqos,                                                      --          .awqos
			m0_awvalid  => h2f_bus_awvalid,                                                    --          .awvalid
			m0_awready  => h2f_bus_awready,                                                    --          .awready
			m0_wdata    => h2f_bus_wdata,                                                      --          .wdata
			m0_wstrb    => h2f_bus_wstrb,                                                      --          .wstrb
			m0_wlast    => h2f_bus_wlast,                                                      --          .wlast
			m0_wvalid   => h2f_bus_wvalid,                                                     --          .wvalid
			m0_wready   => h2f_bus_wready,                                                     --          .wready
			m0_bid      => h2f_bus_bid,                                                        --          .bid
			m0_bresp    => h2f_bus_bresp,                                                      --          .bresp
			m0_bvalid   => h2f_bus_bvalid,                                                     --          .bvalid
			m0_bready   => h2f_bus_bready,                                                     --          .bready
			m0_arid     => h2f_bus_arid,                                                       --          .arid
			m0_araddr   => h2f_bus_araddr,                                                     --          .araddr
			m0_arlen    => h2f_bus_arlen,                                                      --          .arlen
			m0_arsize   => h2f_bus_arsize,                                                     --          .arsize
			m0_arburst  => h2f_bus_arburst,                                                    --          .arburst
			m0_arlock   => h2f_bus_arlock,                                                     --          .arlock
			m0_arcache  => h2f_bus_arcache,                                                    --          .arcache
			m0_arprot   => h2f_bus_arprot,                                                     --          .arprot
			m0_arqos    => h2f_bus_arqos,                                                      --          .arqos
			m0_arvalid  => h2f_bus_arvalid,                                                    --          .arvalid
			m0_arready  => h2f_bus_arready,                                                    --          .arready
			m0_rid      => h2f_bus_rid,                                                        --          .rid
			m0_rdata    => h2f_bus_rdata,                                                      --          .rdata
			m0_rresp    => h2f_bus_rresp,                                                      --          .rresp
			m0_rlast    => h2f_bus_rlast,                                                      --          .rlast
			m0_rvalid   => h2f_bus_rvalid,                                                     --          .rvalid
			m0_rready   => h2f_bus_rready,                                                     --          .rready
			s0_awuser   => "0000000000000000000000000000000000000000000000000000000000000000", -- (terminated)
			s0_awregion => "0000",                                                             -- (terminated)
			s0_wuser    => "0000000000000000000000000000000000000000000000000000000000000000", -- (terminated)
			s0_buser    => open,                                                               -- (terminated)
			s0_aruser   => "0000000000000000000000000000000000000000000000000000000000000000", -- (terminated)
			s0_arregion => "0000",                                                             -- (terminated)
			s0_ruser    => open,                                                               -- (terminated)
			m0_awuser   => open,                                                               -- (terminated)
			m0_awregion => open,                                                               -- (terminated)
			m0_wuser    => open,                                                               -- (terminated)
			m0_buser    => "0000000000000000000000000000000000000000000000000000000000000000", -- (terminated)
			m0_aruser   => open,                                                               -- (terminated)
			m0_arregion => open,                                                               -- (terminated)
			m0_ruser    => "0000000000000000000000000000000000000000000000000000000000000000", -- (terminated)
			m0_wid      => open,                                                               -- (terminated)
			s0_wid      => "000000000000"                                                      -- (terminated)
		);

	buttons_i : component standalone_hps_buttons_i
		port map (
			clk      => clk_clk,                                  --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_1_buttons_i_s1_address,   --                  s1.address
			readdata => mm_interconnect_1_buttons_i_s1_readdata,  --                    .readdata
			in_port  => buttons_i_export                          -- external_connection.export
		);

	dipsw_i : component standalone_hps_buttons_i
		port map (
			clk      => clk_clk,                                  --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_1_dipsw_i_s1_address,     --                  s1.address
			readdata => mm_interconnect_1_dipsw_i_s1_readdata,    --                    .readdata
			in_port  => dipsw_i_export                            -- external_connection.export
		);

	hps_0 : component standalone_hps_hps_0
		generic map (
			F2S_Width => 1,
			S2F_Width => 1
		)
		port map (
			f2h_cold_rst_req_n       => reset_reset_n,                   --  f2h_cold_reset_req.reset_n
			f2h_dbg_rst_req_n        => reset_reset_n,                   -- f2h_debug_reset_req.reset_n
			f2h_warm_rst_req_n       => reset_reset_n,                   --  f2h_warm_reset_req.reset_n
			f2h_stm_hwevents         => open,                            --   f2h_stm_hw_events.stm_hwevents
			mem_a                    => memory_mem_a,                    --              memory.mem_a
			mem_ba                   => memory_mem_ba,                   --                    .mem_ba
			mem_ck                   => memory_mem_ck,                   --                    .mem_ck
			mem_ck_n                 => memory_mem_ck_n,                 --                    .mem_ck_n
			mem_cke                  => memory_mem_cke,                  --                    .mem_cke
			mem_cs_n                 => memory_mem_cs_n,                 --                    .mem_cs_n
			mem_ras_n                => memory_mem_ras_n,                --                    .mem_ras_n
			mem_cas_n                => memory_mem_cas_n,                --                    .mem_cas_n
			mem_we_n                 => memory_mem_we_n,                 --                    .mem_we_n
			mem_reset_n              => memory_mem_reset_n,              --                    .mem_reset_n
			mem_dq                   => memory_mem_dq,                   --                    .mem_dq
			mem_dqs                  => memory_mem_dqs,                  --                    .mem_dqs
			mem_dqs_n                => memory_mem_dqs_n,                --                    .mem_dqs_n
			mem_odt                  => memory_mem_odt,                  --                    .mem_odt
			mem_dm                   => memory_mem_dm,                   --                    .mem_dm
			oct_rzqin                => memory_oct_rzqin,                --                    .oct_rzqin
			hps_io_emac1_inst_TX_CLK => hps_io_hps_io_emac1_inst_TX_CLK, --              hps_io.hps_io_emac1_inst_TX_CLK
			hps_io_emac1_inst_TXD0   => hps_io_hps_io_emac1_inst_TXD0,   --                    .hps_io_emac1_inst_TXD0
			hps_io_emac1_inst_TXD1   => hps_io_hps_io_emac1_inst_TXD1,   --                    .hps_io_emac1_inst_TXD1
			hps_io_emac1_inst_TXD2   => hps_io_hps_io_emac1_inst_TXD2,   --                    .hps_io_emac1_inst_TXD2
			hps_io_emac1_inst_TXD3   => hps_io_hps_io_emac1_inst_TXD3,   --                    .hps_io_emac1_inst_TXD3
			hps_io_emac1_inst_RXD0   => hps_io_hps_io_emac1_inst_RXD0,   --                    .hps_io_emac1_inst_RXD0
			hps_io_emac1_inst_MDIO   => hps_io_hps_io_emac1_inst_MDIO,   --                    .hps_io_emac1_inst_MDIO
			hps_io_emac1_inst_MDC    => hps_io_hps_io_emac1_inst_MDC,    --                    .hps_io_emac1_inst_MDC
			hps_io_emac1_inst_RX_CTL => hps_io_hps_io_emac1_inst_RX_CTL, --                    .hps_io_emac1_inst_RX_CTL
			hps_io_emac1_inst_TX_CTL => hps_io_hps_io_emac1_inst_TX_CTL, --                    .hps_io_emac1_inst_TX_CTL
			hps_io_emac1_inst_RX_CLK => hps_io_hps_io_emac1_inst_RX_CLK, --                    .hps_io_emac1_inst_RX_CLK
			hps_io_emac1_inst_RXD1   => hps_io_hps_io_emac1_inst_RXD1,   --                    .hps_io_emac1_inst_RXD1
			hps_io_emac1_inst_RXD2   => hps_io_hps_io_emac1_inst_RXD2,   --                    .hps_io_emac1_inst_RXD2
			hps_io_emac1_inst_RXD3   => hps_io_hps_io_emac1_inst_RXD3,   --                    .hps_io_emac1_inst_RXD3
			hps_io_qspi_inst_IO0     => hps_io_hps_io_qspi_inst_IO0,     --                    .hps_io_qspi_inst_IO0
			hps_io_qspi_inst_IO1     => hps_io_hps_io_qspi_inst_IO1,     --                    .hps_io_qspi_inst_IO1
			hps_io_qspi_inst_IO2     => hps_io_hps_io_qspi_inst_IO2,     --                    .hps_io_qspi_inst_IO2
			hps_io_qspi_inst_IO3     => hps_io_hps_io_qspi_inst_IO3,     --                    .hps_io_qspi_inst_IO3
			hps_io_qspi_inst_SS0     => hps_io_hps_io_qspi_inst_SS0,     --                    .hps_io_qspi_inst_SS0
			hps_io_qspi_inst_CLK     => hps_io_hps_io_qspi_inst_CLK,     --                    .hps_io_qspi_inst_CLK
			hps_io_sdio_inst_CMD     => hps_io_hps_io_sdio_inst_CMD,     --                    .hps_io_sdio_inst_CMD
			hps_io_sdio_inst_D0      => hps_io_hps_io_sdio_inst_D0,      --                    .hps_io_sdio_inst_D0
			hps_io_sdio_inst_D1      => hps_io_hps_io_sdio_inst_D1,      --                    .hps_io_sdio_inst_D1
			hps_io_sdio_inst_CLK     => hps_io_hps_io_sdio_inst_CLK,     --                    .hps_io_sdio_inst_CLK
			hps_io_sdio_inst_D2      => hps_io_hps_io_sdio_inst_D2,      --                    .hps_io_sdio_inst_D2
			hps_io_sdio_inst_D3      => hps_io_hps_io_sdio_inst_D3,      --                    .hps_io_sdio_inst_D3
			hps_io_usb1_inst_D0      => hps_io_hps_io_usb1_inst_D0,      --                    .hps_io_usb1_inst_D0
			hps_io_usb1_inst_D1      => hps_io_hps_io_usb1_inst_D1,      --                    .hps_io_usb1_inst_D1
			hps_io_usb1_inst_D2      => hps_io_hps_io_usb1_inst_D2,      --                    .hps_io_usb1_inst_D2
			hps_io_usb1_inst_D3      => hps_io_hps_io_usb1_inst_D3,      --                    .hps_io_usb1_inst_D3
			hps_io_usb1_inst_D4      => hps_io_hps_io_usb1_inst_D4,      --                    .hps_io_usb1_inst_D4
			hps_io_usb1_inst_D5      => hps_io_hps_io_usb1_inst_D5,      --                    .hps_io_usb1_inst_D5
			hps_io_usb1_inst_D6      => hps_io_hps_io_usb1_inst_D6,      --                    .hps_io_usb1_inst_D6
			hps_io_usb1_inst_D7      => hps_io_hps_io_usb1_inst_D7,      --                    .hps_io_usb1_inst_D7
			hps_io_usb1_inst_CLK     => hps_io_hps_io_usb1_inst_CLK,     --                    .hps_io_usb1_inst_CLK
			hps_io_usb1_inst_STP     => hps_io_hps_io_usb1_inst_STP,     --                    .hps_io_usb1_inst_STP
			hps_io_usb1_inst_DIR     => hps_io_hps_io_usb1_inst_DIR,     --                    .hps_io_usb1_inst_DIR
			hps_io_usb1_inst_NXT     => hps_io_hps_io_usb1_inst_NXT,     --                    .hps_io_usb1_inst_NXT
			hps_io_spim0_inst_CLK    => hps_io_hps_io_spim0_inst_CLK,    --                    .hps_io_spim0_inst_CLK
			hps_io_spim0_inst_MOSI   => hps_io_hps_io_spim0_inst_MOSI,   --                    .hps_io_spim0_inst_MOSI
			hps_io_spim0_inst_MISO   => hps_io_hps_io_spim0_inst_MISO,   --                    .hps_io_spim0_inst_MISO
			hps_io_spim0_inst_SS0    => hps_io_hps_io_spim0_inst_SS0,    --                    .hps_io_spim0_inst_SS0
			hps_io_uart0_inst_RX     => hps_io_hps_io_uart0_inst_RX,     --                    .hps_io_uart0_inst_RX
			hps_io_uart0_inst_TX     => hps_io_hps_io_uart0_inst_TX,     --                    .hps_io_uart0_inst_TX
			hps_io_i2c0_inst_SDA     => hps_io_hps_io_i2c0_inst_SDA,     --                    .hps_io_i2c0_inst_SDA
			hps_io_i2c0_inst_SCL     => hps_io_hps_io_i2c0_inst_SCL,     --                    .hps_io_i2c0_inst_SCL
			hps_io_can0_inst_RX      => hps_io_hps_io_can0_inst_RX,      --                    .hps_io_can0_inst_RX
			hps_io_can0_inst_TX      => hps_io_hps_io_can0_inst_TX,      --                    .hps_io_can0_inst_TX
			hps_io_trace_inst_CLK    => hps_io_hps_io_trace_inst_CLK,    --                    .hps_io_trace_inst_CLK
			hps_io_trace_inst_D0     => hps_io_hps_io_trace_inst_D0,     --                    .hps_io_trace_inst_D0
			hps_io_trace_inst_D1     => hps_io_hps_io_trace_inst_D1,     --                    .hps_io_trace_inst_D1
			hps_io_trace_inst_D2     => hps_io_hps_io_trace_inst_D2,     --                    .hps_io_trace_inst_D2
			hps_io_trace_inst_D3     => hps_io_hps_io_trace_inst_D3,     --                    .hps_io_trace_inst_D3
			hps_io_trace_inst_D4     => hps_io_hps_io_trace_inst_D4,     --                    .hps_io_trace_inst_D4
			hps_io_trace_inst_D5     => hps_io_hps_io_trace_inst_D5,     --                    .hps_io_trace_inst_D5
			hps_io_trace_inst_D6     => hps_io_hps_io_trace_inst_D6,     --                    .hps_io_trace_inst_D6
			hps_io_trace_inst_D7     => hps_io_hps_io_trace_inst_D7,     --                    .hps_io_trace_inst_D7
			h2f_rst_n                => hps_0_h2f_reset_reset,           --           h2f_reset.reset_n
			h2f_axi_clk              => clk_clk,                         --       h2f_axi_clock.clk
			h2f_AWID                 => hps_0_h2f_axi_master_awid,       --      h2f_axi_master.awid
			h2f_AWADDR               => hps_0_h2f_axi_master_awaddr,     --                    .awaddr
			h2f_AWLEN                => hps_0_h2f_axi_master_awlen,      --                    .awlen
			h2f_AWSIZE               => hps_0_h2f_axi_master_awsize,     --                    .awsize
			h2f_AWBURST              => hps_0_h2f_axi_master_awburst,    --                    .awburst
			h2f_AWLOCK               => hps_0_h2f_axi_master_awlock,     --                    .awlock
			h2f_AWCACHE              => hps_0_h2f_axi_master_awcache,    --                    .awcache
			h2f_AWPROT               => hps_0_h2f_axi_master_awprot,     --                    .awprot
			h2f_AWVALID              => hps_0_h2f_axi_master_awvalid,    --                    .awvalid
			h2f_AWREADY              => hps_0_h2f_axi_master_awready,    --                    .awready
			h2f_WID                  => hps_0_h2f_axi_master_wid,        --                    .wid
			h2f_WDATA                => hps_0_h2f_axi_master_wdata,      --                    .wdata
			h2f_WSTRB                => hps_0_h2f_axi_master_wstrb,      --                    .wstrb
			h2f_WLAST                => hps_0_h2f_axi_master_wlast,      --                    .wlast
			h2f_WVALID               => hps_0_h2f_axi_master_wvalid,     --                    .wvalid
			h2f_WREADY               => hps_0_h2f_axi_master_wready,     --                    .wready
			h2f_BID                  => hps_0_h2f_axi_master_bid,        --                    .bid
			h2f_BRESP                => hps_0_h2f_axi_master_bresp,      --                    .bresp
			h2f_BVALID               => hps_0_h2f_axi_master_bvalid,     --                    .bvalid
			h2f_BREADY               => hps_0_h2f_axi_master_bready,     --                    .bready
			h2f_ARID                 => hps_0_h2f_axi_master_arid,       --                    .arid
			h2f_ARADDR               => hps_0_h2f_axi_master_araddr,     --                    .araddr
			h2f_ARLEN                => hps_0_h2f_axi_master_arlen,      --                    .arlen
			h2f_ARSIZE               => hps_0_h2f_axi_master_arsize,     --                    .arsize
			h2f_ARBURST              => hps_0_h2f_axi_master_arburst,    --                    .arburst
			h2f_ARLOCK               => hps_0_h2f_axi_master_arlock,     --                    .arlock
			h2f_ARCACHE              => hps_0_h2f_axi_master_arcache,    --                    .arcache
			h2f_ARPROT               => hps_0_h2f_axi_master_arprot,     --                    .arprot
			h2f_ARVALID              => hps_0_h2f_axi_master_arvalid,    --                    .arvalid
			h2f_ARREADY              => hps_0_h2f_axi_master_arready,    --                    .arready
			h2f_RID                  => hps_0_h2f_axi_master_rid,        --                    .rid
			h2f_RDATA                => hps_0_h2f_axi_master_rdata,      --                    .rdata
			h2f_RRESP                => hps_0_h2f_axi_master_rresp,      --                    .rresp
			h2f_RLAST                => hps_0_h2f_axi_master_rlast,      --                    .rlast
			h2f_RVALID               => hps_0_h2f_axi_master_rvalid,     --                    .rvalid
			h2f_RREADY               => hps_0_h2f_axi_master_rready,     --                    .rready
			f2h_axi_clk              => clk_clk,                         --       f2h_axi_clock.clk
			f2h_AWID                 => open,                            --       f2h_axi_slave.awid
			f2h_AWADDR               => open,                            --                    .awaddr
			f2h_AWLEN                => open,                            --                    .awlen
			f2h_AWSIZE               => open,                            --                    .awsize
			f2h_AWBURST              => open,                            --                    .awburst
			f2h_AWLOCK               => open,                            --                    .awlock
			f2h_AWCACHE              => open,                            --                    .awcache
			f2h_AWPROT               => open,                            --                    .awprot
			f2h_AWVALID              => open,                            --                    .awvalid
			f2h_AWREADY              => open,                            --                    .awready
			f2h_AWUSER               => open,                            --                    .awuser
			f2h_WID                  => open,                            --                    .wid
			f2h_WDATA                => open,                            --                    .wdata
			f2h_WSTRB                => open,                            --                    .wstrb
			f2h_WLAST                => open,                            --                    .wlast
			f2h_WVALID               => open,                            --                    .wvalid
			f2h_WREADY               => open,                            --                    .wready
			f2h_BID                  => open,                            --                    .bid
			f2h_BRESP                => open,                            --                    .bresp
			f2h_BVALID               => open,                            --                    .bvalid
			f2h_BREADY               => open,                            --                    .bready
			f2h_ARID                 => open,                            --                    .arid
			f2h_ARADDR               => open,                            --                    .araddr
			f2h_ARLEN                => open,                            --                    .arlen
			f2h_ARSIZE               => open,                            --                    .arsize
			f2h_ARBURST              => open,                            --                    .arburst
			f2h_ARLOCK               => open,                            --                    .arlock
			f2h_ARCACHE              => open,                            --                    .arcache
			f2h_ARPROT               => open,                            --                    .arprot
			f2h_ARVALID              => open,                            --                    .arvalid
			f2h_ARREADY              => open,                            --                    .arready
			f2h_ARUSER               => open,                            --                    .aruser
			f2h_RID                  => open,                            --                    .rid
			f2h_RDATA                => open,                            --                    .rdata
			f2h_RRESP                => open,                            --                    .rresp
			f2h_RLAST                => open,                            --                    .rlast
			f2h_RVALID               => open,                            --                    .rvalid
			f2h_RREADY               => open,                            --                    .rready
			h2f_lw_axi_clk           => clk_clk,                         --    h2f_lw_axi_clock.clk
			h2f_lw_AWID              => hps_0_h2f_lw_axi_master_awid,    --   h2f_lw_axi_master.awid
			h2f_lw_AWADDR            => hps_0_h2f_lw_axi_master_awaddr,  --                    .awaddr
			h2f_lw_AWLEN             => hps_0_h2f_lw_axi_master_awlen,   --                    .awlen
			h2f_lw_AWSIZE            => hps_0_h2f_lw_axi_master_awsize,  --                    .awsize
			h2f_lw_AWBURST           => hps_0_h2f_lw_axi_master_awburst, --                    .awburst
			h2f_lw_AWLOCK            => hps_0_h2f_lw_axi_master_awlock,  --                    .awlock
			h2f_lw_AWCACHE           => hps_0_h2f_lw_axi_master_awcache, --                    .awcache
			h2f_lw_AWPROT            => hps_0_h2f_lw_axi_master_awprot,  --                    .awprot
			h2f_lw_AWVALID           => hps_0_h2f_lw_axi_master_awvalid, --                    .awvalid
			h2f_lw_AWREADY           => hps_0_h2f_lw_axi_master_awready, --                    .awready
			h2f_lw_WID               => hps_0_h2f_lw_axi_master_wid,     --                    .wid
			h2f_lw_WDATA             => hps_0_h2f_lw_axi_master_wdata,   --                    .wdata
			h2f_lw_WSTRB             => hps_0_h2f_lw_axi_master_wstrb,   --                    .wstrb
			h2f_lw_WLAST             => hps_0_h2f_lw_axi_master_wlast,   --                    .wlast
			h2f_lw_WVALID            => hps_0_h2f_lw_axi_master_wvalid,  --                    .wvalid
			h2f_lw_WREADY            => hps_0_h2f_lw_axi_master_wready,  --                    .wready
			h2f_lw_BID               => hps_0_h2f_lw_axi_master_bid,     --                    .bid
			h2f_lw_BRESP             => hps_0_h2f_lw_axi_master_bresp,   --                    .bresp
			h2f_lw_BVALID            => hps_0_h2f_lw_axi_master_bvalid,  --                    .bvalid
			h2f_lw_BREADY            => hps_0_h2f_lw_axi_master_bready,  --                    .bready
			h2f_lw_ARID              => hps_0_h2f_lw_axi_master_arid,    --                    .arid
			h2f_lw_ARADDR            => hps_0_h2f_lw_axi_master_araddr,  --                    .araddr
			h2f_lw_ARLEN             => hps_0_h2f_lw_axi_master_arlen,   --                    .arlen
			h2f_lw_ARSIZE            => hps_0_h2f_lw_axi_master_arsize,  --                    .arsize
			h2f_lw_ARBURST           => hps_0_h2f_lw_axi_master_arburst, --                    .arburst
			h2f_lw_ARLOCK            => hps_0_h2f_lw_axi_master_arlock,  --                    .arlock
			h2f_lw_ARCACHE           => hps_0_h2f_lw_axi_master_arcache, --                    .arcache
			h2f_lw_ARPROT            => hps_0_h2f_lw_axi_master_arprot,  --                    .arprot
			h2f_lw_ARVALID           => hps_0_h2f_lw_axi_master_arvalid, --                    .arvalid
			h2f_lw_ARREADY           => hps_0_h2f_lw_axi_master_arready, --                    .arready
			h2f_lw_RID               => hps_0_h2f_lw_axi_master_rid,     --                    .rid
			h2f_lw_RDATA             => hps_0_h2f_lw_axi_master_rdata,   --                    .rdata
			h2f_lw_RRESP             => hps_0_h2f_lw_axi_master_rresp,   --                    .rresp
			h2f_lw_RLAST             => hps_0_h2f_lw_axi_master_rlast,   --                    .rlast
			h2f_lw_RVALID            => hps_0_h2f_lw_axi_master_rvalid,  --                    .rvalid
			h2f_lw_RREADY            => hps_0_h2f_lw_axi_master_rready,  --                    .rready
			f2h_irq_p0               => hps_0_f2h_irq0_irq,              --            f2h_irq0.irq
			f2h_irq_p1               => hps_0_f2h_irq1_irq               --            f2h_irq1.irq
		);

	leds_o : component standalone_hps_leds_o
		port map (
			clk        => clk_clk,                                     --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,    --               reset.reset_n
			address    => mm_interconnect_1_leds_o_s1_address,         --                  s1.address
			write_n    => mm_interconnect_1_leds_o_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_1_leds_o_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_1_leds_o_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_1_leds_o_s1_readdata,        --                    .readdata
			out_port   => leds_o_export                                -- external_connection.export
		);

	mm_interconnect_0 : component standalone_hps_mm_interconnect_0
		port map (
			axi_bridge_0_s0_awid                               => mm_interconnect_0_axi_bridge_0_s0_awid,    --                              axi_bridge_0_s0.awid
			axi_bridge_0_s0_awaddr                             => mm_interconnect_0_axi_bridge_0_s0_awaddr,  --                                             .awaddr
			axi_bridge_0_s0_awlen                              => mm_interconnect_0_axi_bridge_0_s0_awlen,   --                                             .awlen
			axi_bridge_0_s0_awsize                             => mm_interconnect_0_axi_bridge_0_s0_awsize,  --                                             .awsize
			axi_bridge_0_s0_awburst                            => mm_interconnect_0_axi_bridge_0_s0_awburst, --                                             .awburst
			axi_bridge_0_s0_awlock                             => mm_interconnect_0_axi_bridge_0_s0_awlock,  --                                             .awlock
			axi_bridge_0_s0_awcache                            => mm_interconnect_0_axi_bridge_0_s0_awcache, --                                             .awcache
			axi_bridge_0_s0_awprot                             => mm_interconnect_0_axi_bridge_0_s0_awprot,  --                                             .awprot
			axi_bridge_0_s0_awqos                              => mm_interconnect_0_axi_bridge_0_s0_awqos,   --                                             .awqos
			axi_bridge_0_s0_awvalid                            => mm_interconnect_0_axi_bridge_0_s0_awvalid, --                                             .awvalid
			axi_bridge_0_s0_awready                            => mm_interconnect_0_axi_bridge_0_s0_awready, --                                             .awready
			axi_bridge_0_s0_wdata                              => mm_interconnect_0_axi_bridge_0_s0_wdata,   --                                             .wdata
			axi_bridge_0_s0_wstrb                              => mm_interconnect_0_axi_bridge_0_s0_wstrb,   --                                             .wstrb
			axi_bridge_0_s0_wlast                              => mm_interconnect_0_axi_bridge_0_s0_wlast,   --                                             .wlast
			axi_bridge_0_s0_wvalid                             => mm_interconnect_0_axi_bridge_0_s0_wvalid,  --                                             .wvalid
			axi_bridge_0_s0_wready                             => mm_interconnect_0_axi_bridge_0_s0_wready,  --                                             .wready
			axi_bridge_0_s0_bid                                => mm_interconnect_0_axi_bridge_0_s0_bid,     --                                             .bid
			axi_bridge_0_s0_bresp                              => mm_interconnect_0_axi_bridge_0_s0_bresp,   --                                             .bresp
			axi_bridge_0_s0_bvalid                             => mm_interconnect_0_axi_bridge_0_s0_bvalid,  --                                             .bvalid
			axi_bridge_0_s0_bready                             => mm_interconnect_0_axi_bridge_0_s0_bready,  --                                             .bready
			axi_bridge_0_s0_arid                               => mm_interconnect_0_axi_bridge_0_s0_arid,    --                                             .arid
			axi_bridge_0_s0_araddr                             => mm_interconnect_0_axi_bridge_0_s0_araddr,  --                                             .araddr
			axi_bridge_0_s0_arlen                              => mm_interconnect_0_axi_bridge_0_s0_arlen,   --                                             .arlen
			axi_bridge_0_s0_arsize                             => mm_interconnect_0_axi_bridge_0_s0_arsize,  --                                             .arsize
			axi_bridge_0_s0_arburst                            => mm_interconnect_0_axi_bridge_0_s0_arburst, --                                             .arburst
			axi_bridge_0_s0_arlock                             => mm_interconnect_0_axi_bridge_0_s0_arlock,  --                                             .arlock
			axi_bridge_0_s0_arcache                            => mm_interconnect_0_axi_bridge_0_s0_arcache, --                                             .arcache
			axi_bridge_0_s0_arprot                             => mm_interconnect_0_axi_bridge_0_s0_arprot,  --                                             .arprot
			axi_bridge_0_s0_arqos                              => mm_interconnect_0_axi_bridge_0_s0_arqos,   --                                             .arqos
			axi_bridge_0_s0_arvalid                            => mm_interconnect_0_axi_bridge_0_s0_arvalid, --                                             .arvalid
			axi_bridge_0_s0_arready                            => mm_interconnect_0_axi_bridge_0_s0_arready, --                                             .arready
			axi_bridge_0_s0_rid                                => mm_interconnect_0_axi_bridge_0_s0_rid,     --                                             .rid
			axi_bridge_0_s0_rdata                              => mm_interconnect_0_axi_bridge_0_s0_rdata,   --                                             .rdata
			axi_bridge_0_s0_rresp                              => mm_interconnect_0_axi_bridge_0_s0_rresp,   --                                             .rresp
			axi_bridge_0_s0_rlast                              => mm_interconnect_0_axi_bridge_0_s0_rlast,   --                                             .rlast
			axi_bridge_0_s0_rvalid                             => mm_interconnect_0_axi_bridge_0_s0_rvalid,  --                                             .rvalid
			axi_bridge_0_s0_rready                             => mm_interconnect_0_axi_bridge_0_s0_rready,  --                                             .rready
			hps_0_h2f_axi_master_awid                          => hps_0_h2f_axi_master_awid,                 --                         hps_0_h2f_axi_master.awid
			hps_0_h2f_axi_master_awaddr                        => hps_0_h2f_axi_master_awaddr,               --                                             .awaddr
			hps_0_h2f_axi_master_awlen                         => hps_0_h2f_axi_master_awlen,                --                                             .awlen
			hps_0_h2f_axi_master_awsize                        => hps_0_h2f_axi_master_awsize,               --                                             .awsize
			hps_0_h2f_axi_master_awburst                       => hps_0_h2f_axi_master_awburst,              --                                             .awburst
			hps_0_h2f_axi_master_awlock                        => hps_0_h2f_axi_master_awlock,               --                                             .awlock
			hps_0_h2f_axi_master_awcache                       => hps_0_h2f_axi_master_awcache,              --                                             .awcache
			hps_0_h2f_axi_master_awprot                        => hps_0_h2f_axi_master_awprot,               --                                             .awprot
			hps_0_h2f_axi_master_awvalid                       => hps_0_h2f_axi_master_awvalid,              --                                             .awvalid
			hps_0_h2f_axi_master_awready                       => hps_0_h2f_axi_master_awready,              --                                             .awready
			hps_0_h2f_axi_master_wid                           => hps_0_h2f_axi_master_wid,                  --                                             .wid
			hps_0_h2f_axi_master_wdata                         => hps_0_h2f_axi_master_wdata,                --                                             .wdata
			hps_0_h2f_axi_master_wstrb                         => hps_0_h2f_axi_master_wstrb,                --                                             .wstrb
			hps_0_h2f_axi_master_wlast                         => hps_0_h2f_axi_master_wlast,                --                                             .wlast
			hps_0_h2f_axi_master_wvalid                        => hps_0_h2f_axi_master_wvalid,               --                                             .wvalid
			hps_0_h2f_axi_master_wready                        => hps_0_h2f_axi_master_wready,               --                                             .wready
			hps_0_h2f_axi_master_bid                           => hps_0_h2f_axi_master_bid,                  --                                             .bid
			hps_0_h2f_axi_master_bresp                         => hps_0_h2f_axi_master_bresp,                --                                             .bresp
			hps_0_h2f_axi_master_bvalid                        => hps_0_h2f_axi_master_bvalid,               --                                             .bvalid
			hps_0_h2f_axi_master_bready                        => hps_0_h2f_axi_master_bready,               --                                             .bready
			hps_0_h2f_axi_master_arid                          => hps_0_h2f_axi_master_arid,                 --                                             .arid
			hps_0_h2f_axi_master_araddr                        => hps_0_h2f_axi_master_araddr,               --                                             .araddr
			hps_0_h2f_axi_master_arlen                         => hps_0_h2f_axi_master_arlen,                --                                             .arlen
			hps_0_h2f_axi_master_arsize                        => hps_0_h2f_axi_master_arsize,               --                                             .arsize
			hps_0_h2f_axi_master_arburst                       => hps_0_h2f_axi_master_arburst,              --                                             .arburst
			hps_0_h2f_axi_master_arlock                        => hps_0_h2f_axi_master_arlock,               --                                             .arlock
			hps_0_h2f_axi_master_arcache                       => hps_0_h2f_axi_master_arcache,              --                                             .arcache
			hps_0_h2f_axi_master_arprot                        => hps_0_h2f_axi_master_arprot,               --                                             .arprot
			hps_0_h2f_axi_master_arvalid                       => hps_0_h2f_axi_master_arvalid,              --                                             .arvalid
			hps_0_h2f_axi_master_arready                       => hps_0_h2f_axi_master_arready,              --                                             .arready
			hps_0_h2f_axi_master_rid                           => hps_0_h2f_axi_master_rid,                  --                                             .rid
			hps_0_h2f_axi_master_rdata                         => hps_0_h2f_axi_master_rdata,                --                                             .rdata
			hps_0_h2f_axi_master_rresp                         => hps_0_h2f_axi_master_rresp,                --                                             .rresp
			hps_0_h2f_axi_master_rlast                         => hps_0_h2f_axi_master_rlast,                --                                             .rlast
			hps_0_h2f_axi_master_rvalid                        => hps_0_h2f_axi_master_rvalid,               --                                             .rvalid
			hps_0_h2f_axi_master_rready                        => hps_0_h2f_axi_master_rready,               --                                             .rready
			clk_0_clk_clk                                      => clk_clk,                                   --                                    clk_0_clk.clk
			axi_bridge_0_clk_reset_reset_bridge_in_reset_reset => rst_controller_reset_out_reset             -- axi_bridge_0_clk_reset_reset_bridge_in_reset.reset
		);

	mm_interconnect_1 : component standalone_hps_mm_interconnect_1
		port map (
			hps_0_h2f_lw_axi_master_awid                                        => hps_0_h2f_lw_axi_master_awid,            --                                       hps_0_h2f_lw_axi_master.awid
			hps_0_h2f_lw_axi_master_awaddr                                      => hps_0_h2f_lw_axi_master_awaddr,          --                                                              .awaddr
			hps_0_h2f_lw_axi_master_awlen                                       => hps_0_h2f_lw_axi_master_awlen,           --                                                              .awlen
			hps_0_h2f_lw_axi_master_awsize                                      => hps_0_h2f_lw_axi_master_awsize,          --                                                              .awsize
			hps_0_h2f_lw_axi_master_awburst                                     => hps_0_h2f_lw_axi_master_awburst,         --                                                              .awburst
			hps_0_h2f_lw_axi_master_awlock                                      => hps_0_h2f_lw_axi_master_awlock,          --                                                              .awlock
			hps_0_h2f_lw_axi_master_awcache                                     => hps_0_h2f_lw_axi_master_awcache,         --                                                              .awcache
			hps_0_h2f_lw_axi_master_awprot                                      => hps_0_h2f_lw_axi_master_awprot,          --                                                              .awprot
			hps_0_h2f_lw_axi_master_awvalid                                     => hps_0_h2f_lw_axi_master_awvalid,         --                                                              .awvalid
			hps_0_h2f_lw_axi_master_awready                                     => hps_0_h2f_lw_axi_master_awready,         --                                                              .awready
			hps_0_h2f_lw_axi_master_wid                                         => hps_0_h2f_lw_axi_master_wid,             --                                                              .wid
			hps_0_h2f_lw_axi_master_wdata                                       => hps_0_h2f_lw_axi_master_wdata,           --                                                              .wdata
			hps_0_h2f_lw_axi_master_wstrb                                       => hps_0_h2f_lw_axi_master_wstrb,           --                                                              .wstrb
			hps_0_h2f_lw_axi_master_wlast                                       => hps_0_h2f_lw_axi_master_wlast,           --                                                              .wlast
			hps_0_h2f_lw_axi_master_wvalid                                      => hps_0_h2f_lw_axi_master_wvalid,          --                                                              .wvalid
			hps_0_h2f_lw_axi_master_wready                                      => hps_0_h2f_lw_axi_master_wready,          --                                                              .wready
			hps_0_h2f_lw_axi_master_bid                                         => hps_0_h2f_lw_axi_master_bid,             --                                                              .bid
			hps_0_h2f_lw_axi_master_bresp                                       => hps_0_h2f_lw_axi_master_bresp,           --                                                              .bresp
			hps_0_h2f_lw_axi_master_bvalid                                      => hps_0_h2f_lw_axi_master_bvalid,          --                                                              .bvalid
			hps_0_h2f_lw_axi_master_bready                                      => hps_0_h2f_lw_axi_master_bready,          --                                                              .bready
			hps_0_h2f_lw_axi_master_arid                                        => hps_0_h2f_lw_axi_master_arid,            --                                                              .arid
			hps_0_h2f_lw_axi_master_araddr                                      => hps_0_h2f_lw_axi_master_araddr,          --                                                              .araddr
			hps_0_h2f_lw_axi_master_arlen                                       => hps_0_h2f_lw_axi_master_arlen,           --                                                              .arlen
			hps_0_h2f_lw_axi_master_arsize                                      => hps_0_h2f_lw_axi_master_arsize,          --                                                              .arsize
			hps_0_h2f_lw_axi_master_arburst                                     => hps_0_h2f_lw_axi_master_arburst,         --                                                              .arburst
			hps_0_h2f_lw_axi_master_arlock                                      => hps_0_h2f_lw_axi_master_arlock,          --                                                              .arlock
			hps_0_h2f_lw_axi_master_arcache                                     => hps_0_h2f_lw_axi_master_arcache,         --                                                              .arcache
			hps_0_h2f_lw_axi_master_arprot                                      => hps_0_h2f_lw_axi_master_arprot,          --                                                              .arprot
			hps_0_h2f_lw_axi_master_arvalid                                     => hps_0_h2f_lw_axi_master_arvalid,         --                                                              .arvalid
			hps_0_h2f_lw_axi_master_arready                                     => hps_0_h2f_lw_axi_master_arready,         --                                                              .arready
			hps_0_h2f_lw_axi_master_rid                                         => hps_0_h2f_lw_axi_master_rid,             --                                                              .rid
			hps_0_h2f_lw_axi_master_rdata                                       => hps_0_h2f_lw_axi_master_rdata,           --                                                              .rdata
			hps_0_h2f_lw_axi_master_rresp                                       => hps_0_h2f_lw_axi_master_rresp,           --                                                              .rresp
			hps_0_h2f_lw_axi_master_rlast                                       => hps_0_h2f_lw_axi_master_rlast,           --                                                              .rlast
			hps_0_h2f_lw_axi_master_rvalid                                      => hps_0_h2f_lw_axi_master_rvalid,          --                                                              .rvalid
			hps_0_h2f_lw_axi_master_rready                                      => hps_0_h2f_lw_axi_master_rready,          --                                                              .rready
			clk_0_clk_clk                                                       => clk_clk,                                 --                                                     clk_0_clk.clk
			hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset => rst_controller_001_reset_out_reset,      -- hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
			leds_o_reset_reset_bridge_in_reset_reset                            => rst_controller_reset_out_reset,          --                            leds_o_reset_reset_bridge_in_reset.reset
			buttons_i_s1_address                                                => mm_interconnect_1_buttons_i_s1_address,  --                                                  buttons_i_s1.address
			buttons_i_s1_readdata                                               => mm_interconnect_1_buttons_i_s1_readdata, --                                                              .readdata
			dipsw_i_s1_address                                                  => mm_interconnect_1_dipsw_i_s1_address,    --                                                    dipsw_i_s1.address
			dipsw_i_s1_readdata                                                 => mm_interconnect_1_dipsw_i_s1_readdata,   --                                                              .readdata
			leds_o_s1_address                                                   => mm_interconnect_1_leds_o_s1_address,     --                                                     leds_o_s1.address
			leds_o_s1_write                                                     => mm_interconnect_1_leds_o_s1_write,       --                                                              .write
			leds_o_s1_readdata                                                  => mm_interconnect_1_leds_o_s1_readdata,    --                                                              .readdata
			leds_o_s1_writedata                                                 => mm_interconnect_1_leds_o_s1_writedata,   --                                                              .writedata
			leds_o_s1_chipselect                                                => mm_interconnect_1_leds_o_s1_chipselect   --                                                              .chipselect
		);

	irq_mapper : component standalone_hps_irq_mapper
		port map (
			clk        => open,               --       clk.clk
			reset      => open,               -- clk_reset.reset
			sender_irq => hps_0_f2h_irq0_irq  --    sender.irq
		);

	irq_mapper_001 : component standalone_hps_irq_mapper
		port map (
			clk        => open,               --       clk.clk
			reset      => open,               -- clk_reset.reset
			sender_irq => hps_0_f2h_irq1_irq  --    sender.irq
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,        -- reset_in0.reset
			clk            => clk_clk,                        --       clk.clk
			reset_out      => rst_controller_reset_out_reset, -- reset_out.reset
			reset_req      => open,                           -- (terminated)
			reset_req_in0  => '0',                            -- (terminated)
			reset_in1      => '0',                            -- (terminated)
			reset_req_in1  => '0',                            -- (terminated)
			reset_in2      => '0',                            -- (terminated)
			reset_req_in2  => '0',                            -- (terminated)
			reset_in3      => '0',                            -- (terminated)
			reset_req_in3  => '0',                            -- (terminated)
			reset_in4      => '0',                            -- (terminated)
			reset_req_in4  => '0',                            -- (terminated)
			reset_in5      => '0',                            -- (terminated)
			reset_req_in5  => '0',                            -- (terminated)
			reset_in6      => '0',                            -- (terminated)
			reset_req_in6  => '0',                            -- (terminated)
			reset_in7      => '0',                            -- (terminated)
			reset_req_in7  => '0',                            -- (terminated)
			reset_in8      => '0',                            -- (terminated)
			reset_req_in8  => '0',                            -- (terminated)
			reset_in9      => '0',                            -- (terminated)
			reset_req_in9  => '0',                            -- (terminated)
			reset_in10     => '0',                            -- (terminated)
			reset_req_in10 => '0',                            -- (terminated)
			reset_in11     => '0',                            -- (terminated)
			reset_req_in11 => '0',                            -- (terminated)
			reset_in12     => '0',                            -- (terminated)
			reset_req_in12 => '0',                            -- (terminated)
			reset_in13     => '0',                            -- (terminated)
			reset_req_in13 => '0',                            -- (terminated)
			reset_in14     => '0',                            -- (terminated)
			reset_req_in14 => '0',                            -- (terminated)
			reset_in15     => '0',                            -- (terminated)
			reset_req_in15 => '0'                             -- (terminated)
		);

	rst_controller_001 : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => h2f_reset_reset_n_ports_inv,        -- reset_in0.reset
			clk            => clk_clk,                            --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	h2f_reset_reset_n_ports_inv <= not hps_0_h2f_reset_reset;

	reset_reset_n_ports_inv <= not reset_reset_n;

	mm_interconnect_1_leds_o_s1_write_ports_inv <= not mm_interconnect_1_leds_o_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

	h2f_reset_reset_n <= hps_0_h2f_reset_reset;

end architecture rtl; -- of standalone_hps
