// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 01:35:05 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
WRQLeTfb12ZZGAv5DFAnT9CrP6tOT7x097m6nBiIOmk0v/Y4/aSNopF6ZeAuBmO3
iLYIBWd5CoLuCVWrZqscvTLyTVF9zMBYe1xkMh51/15j7rzcjPIQgUE6ZvMAM3EZ
xXCmuI2dZmEdDUplUHpAUdmTAz1YBkgYUwshLLvOxuA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 32640)
Hfk8S5KmSj1WIINOEMXeAgdf+w1VcG3DMFJEH1CAJg2YeE2ko0rwNCIilJHy5LI8
rJfyxc0W5+b9VkL4HCZf51OwOoBl2KZfn4DVNCBSCbx4g/BcYrGmyqrxM/3a4OEu
zers532raNXZIcVuSW8mohW+mQ9G88kCY+aVi83QJDDUueetyJxB31wbehVCN+1V
Lh53Nhb9v3TrYtnZto7HmEBghFABIRfzYRaOpTREVkRFCPMameOHjJzTWmnYS9Vk
ycDEBXwIZeXznSeMPxma2M1W6he5uunrXXjjfgW7yW2B7rTMbsY1DcCVcJOUBoft
eQk9eeH4w+4ups+aXkzzp9zY5xyZ7l+K0kxiWjRV5ELYALl+NrQqiYSx0Wkrz8br
XbWXbA5i71/vrONDIX2Rz/A6/4UXVJ98Kg5sJ7ajphRL0sqfplRv+tkwNBNxjK0R
GhihnIWkRbpijj40N4GsoFIc/OkfUBvv2A9LA4wMr3cOJT8nEn6yZEOHes/s0a91
CSCT6qfWDYwi1O2e1wG6UNa7y286fxmyrqN1rfa2W+o8LNQ5bd4AYin2XFD2fypa
JC/N9lg3dU0cgh8khkYbGhabIjxb1ngggR+QAVWfbrwVyS7MNqp+AYcu/KSe/9hk
Y1mQ4zRjJXKjXfCg0jhRJJN3kyaalklk5wkBhZ4BoCoT3xn9TYtjfQGzax8b5sDV
ODSV6sen029LyOUr/6G7wqIwqOAwngPUxSkQQ83RRTzT/llNgdgKNynVdYoO+p3m
l7PsOcFxe0iPLvrkZR0Ne4zFbLl1g6oMW1XjNHN0KCqkwW3v+jKFCIRySuOyeC3s
L8fL+TtGjQqOvpL1ZcFFzXx0g62VtBDAzV5hbEUS8NSVB/wl5WeVTFsV/lV04gm9
qQpIhU8Xdnaq3WmbLuabN01euW5vMlNR8bZ4yr/dEKFZ+qYkpOb2UQ29EXmNN5H+
r5N8NRcnex5bmr35M4Fsoux5KtgBKQwFIesL4CzE3Ee+nI3V26G6sfB6Ds4cdXwr
i+C/IibvwN1igAgLJETymSbx1xey+FR5y8bakmXVx4x6tT9QP6/EIOPzH3LrQs6I
7dybmOKK9z5DboVc2BtVw6jEzXDauo5BLBVPe4uyEi9Klqla3uZd2yMzoP/pdwIl
bgQ5VVNWQg8Yq2dhv2gZ0YLw9kabFzSnTc6VDJdM+bPRbfr5eXk+wXvDiRs9xedD
Vncv3QtZS5IBPueLrSs95sfR2S9TRMHg+rQcOUEhekwHCyFUbLj7PElAKEii4VLy
XTOEqrM98X5E2BXGuj2KyuvrsPgA/tqmvQ03f/Iu9W3f6ScJdeb6/QSNBOquHvLw
Fumz5BMYz2N3SNFd8PQ4Bj5rTEVE/NnWTrSnGMVbZPdR73bw4nNJFkAUDSp+D6qO
TyODEEs3D04rotTf3msA3IovhAFSdM1pEMoDl/Z47PipI7MdzZeJy3IEZ10MzLzV
gw8xwhbU7tNlJsFw1DMfy58RYZ5g4iGo8YJieisvJKktiFW7Dj+ueMnu9ZQU5dnw
iDc2jPLKWNiXJo269fobHNf7t6dHR2se3meDNuYJWdg7L8lzFtv/ZBFAhvrNLvUY
NUNr1yjFAJOCS5fQnml1h8Bbfrc+64637O0wAf9SsEBLS99Q3xnrOI2y5vEIdEKL
Ahdy1t7Mr2rOi6spnMShu9ngMH5NoxfUZTe4EZu6X2GNaSOORWbB4AFMucg+N4YU
v5xV//1xGZkUT1BHrQEd4llACgx8tmdBD2OtzBvyc+sDPHYMAYrvKzfxcGOCeYr5
N+B/rhtlFfdQrJnUp1wtqZ+bMivOj+D1SfmxbBbjpP7NGj+NcTTeIve5kQwzOAPZ
bslPO20QLuwa02lBMZaANJuAZZ6CBuSd3pp1QJroHQMzaOsQm3Yk5sX7/IksHgij
2L3i15d35p8NTr/fQdyHsyBaRcKs8hU9ZGR08kt1/J7yneT1JauljS/EG5F1zlg0
t//MsB8lDiVdfXW3KyKdPbh6w0TGUWWzJyiL8IDFB2dwmgcnolID9Y8aaWZJN2Zy
NrUwBYhAqjyURM8h2NhXt+ylMU1PZ3qb51TFDU1l8UcwP43RKEfE792fB/myr2IP
JkPmCnoUsIu2y6tkBK7cIXtM8AtvaE/kn35GMm6vxTSXfzOnRIO8Ih4kwfTAh9EV
51V2srDJobzoS6lWAH1BZ2K09cwNFrpIGpMANM0m9wuwicLQNfat5Xhxk1szJNdD
xrO4ukxjCT7u03GCh9dubZo3n8kKe9QQi34aSeUt56LynF/ESFcoA2xd27brRiW3
UI2E75Wn/X0xdEY8jKEUmIjUxLgBeO2eObo089L9MhBfoD+jvSGmwmmcKqqZowxO
i2Nd1zzsO2KpqjFPCUUizZy1hrmaZeS7RNBBL41vSCzMs2RVAA1VqmfGJPmlsqAJ
XO0udwJNuPxcDabb7EBxewqmMuf4eqEwWfTu9i/aURWTLtZwpyMQvKHR5E15mAyi
yqXCQLaM6fgSThxYQvjHLQZYBCPXaIOI62CUnENdOdkwSUMWYTzzIDgVJ0EYJ4Lp
ePygR72f4mjsS+5IVqH/l4rjs1ioPC7ep70hHHnsKyFJJny3ANTyne3cO+5I0fQ7
yveM6vZczWaGnYlDKUN+pUGbxpSdPzt+iyfeppAO8oBP6MAGbdW8tzFVhvHEC7+X
5bd9NwohnKu8u5qpHBkemd4GbcvNlIcVi9/bEELY+AAibniTHAkKS50chSMaVW2s
CEZTfnQDQ40+ByCbih8VbLOSByxaD9m1QB1OQ05i4LAFZfHTBlUcEu4k559rahRY
T8piSoYrHSXm95bH5Z5CJyzpegAJR3ZSpIxuTvSMRh2ocBA+D+5j+Hljg1afWZSa
43RXi4wCmMB8MwF3N8OYr1ni08ARX739SdIkycl11b8K2rUF6ABK81YKI+EaIHRM
Jv20EpzmI0hDJmRA4Ish38lpWq/nKTLYJC9s7cm80hSWtlxk7tT5LBcnlS7/Sjp2
MC2trRuf+vb98Y0HGcAdZeO4gUMLN8reUyAxnKWJWLTGL5PwO5+/j2ZbUTHy34He
iN/HOiHsWeHhRq4SXAr2oWBw3D8v4OiNhB8MbiA8oiI4dqaiMjzpYOWCElsdMpaF
gEf7iSadtOFoMlbFiEZQlKkfuacgSsrhT8DPavM44c0hitpasSNPlLi1INbqlxe7
amLJ+sL5yDBwOzcY8jt8vVS0lxdxH73qdDoIFkl5rqhPSUSrqUEH6YPqM59AzxMf
NOFo9HCfHQp5TvZXTO2gX0ymRcuR/TVxDpMW5I6Dh2bOrjZIUV4qxCURjyU0px14
+Kl1dZYT/RHl03h94qBInELfsaaQ5xS5tc6bqP84iJLa2XJXXSAL4gl53lakUP0W
CViLm2kE9BNjfhlSJgxHQYAmDJuzcpUHvJBNUyzqMab5A9SI61YVMXSS7EvN4CTE
fNH1QaZrk5Q67My7/3ipbPUB/WrbTi+68dfudgawP8VDRll31fPc+/vV29gczCIz
4pe8XI/CRUwhRtYIUhbZBpkudhPjJYPkGav0IMmEqspagqtBmTWRuNDiXRKFLDuH
HXYxegGap8HVHBDhL4yes4r1FYogRPGv5jl+yJU2zdB/D6tA5fl10Fk9oKrQDCaP
WmZCklzv/Ux1a1LJlpXgaZ8wSrN3+VigVd47/IwE5uTqyQrBFSfZPXZncoNHDiXu
GalZR2cNpTxWAH/9x+avgD0eLe0wL4AXpBdgRCnyPovdz6A0sNXlz+0LOU18ads1
W+nbt1MnZ0Hfn8f767Ph7DMUF9ra8eu6/vSXBYHC8Pr+VqQV9NeOH4RJX+JZZX80
+DUcTR+aCQNbSyzcxGRsqdVlZTQnmaEES6kpSKTt6BodJhr1117z2e7886zFdWtT
TOtUMPf9Ku+5LV2fu/BrP5U19D/S2wOIpobzqgOcQDEc/0id/8ILKnK5BNMJ/bGL
pdRf5lMiJU8LpZq6WoLh61Px+3H1Cx1w6ISfx2/LrdtjrRueIrZp636mikf65s7k
EV2W6C/12fcp2d+jgwL/fXYCMQLWSSq6+4KH/HkI96hUbcoQTGEjNkHDT2idXNFF
JBNwn+l8yF8iA4fQGc8dm9sLdMBIickRsB7uMPBQSJnBDti2j2j/Kg8LPhUkVYYk
cKc/rgrly6IAObfR8uYc+JxrAOoPUXakxcu/lQWRG8q5YQde4ojuyYb9wBgXrVob
JiYx9dPQ/WfOesIUb1VCu5lMVNjBRhOi7sX4m6KcYZDyIP3H2YZ9P5hSrdhLksLF
MGd5HXCuC6t7mffZHXah0z9nx1Dd7EzktS46INXnsognAf/j7zW3R3kllfTWEOyw
pFT/s7q0m1zkZboXXTASuEpRCaTZ3/Fuk0Es0EICtw8zGIMQ9CjHuL0NwOhIkIty
q1G4UpjCqBAgxGTaOQDSRvXmJNzpSGpQgTRI49q1+K0XHHx/LcFkL4RdyF4xh54s
k1lgblwghxsgu9zJQfiVfFNufGmYmf0i9aAMz7J3FylZu0qQg9fnZYG0hYPv7TwB
bvJ4nbco5SsegIEKdGycoURKgjf0LkAFVd9RcOQqR5kxD5BX28KBUGh5zQwbhvkn
Cj4eEnkJGBZ7ZOZDlBoV+mjr+qq0183yWFTxVLi65dFGRgOlNlEruV6v703d9cXM
++e5KQuS5LAW/D1hacAJkIxb0FbQ6bo+2oq+dKDaABXceQRVywW1Y2D8tOOfL/TG
4OMrDN/r0mInpfBeoNeZgBdQr+ReOFQsAXHaIn46GxSMLrxHbgppaQ97/UKsf+Zg
WDaSKRL6FKjmgtYL9uhUQSW7IUPb0RM0+IBmrheudWVz45JxjWewbzJx3Ur0UPt0
3SjhI3U0HfKUBJ0CTela6mdbNOYFi/ONfOfx2UT0SMigj0fp9QcATSNr4zI2/Lo5
BDgkKa2FMRiKUB5FT2QzjS4zg8Cw4gaMTeqKmV1vxCALWyqZr84O5bqmMPh78NCa
Pt0f3/A7EKDF+rCt+F78hd0y9nttCppHk/LHD1fc2k9BNsYNDaM24m4fqLguDx9q
ACCo6O+gZVg4VvUX7AuUw+JN4kwoMUqsrwwjBotccw798RC+Va/3i68JvVUlSMLb
RCuZLnta2XKCrVio1YKJkV0Ku/pKG9fWJQkXDAbvZZPVj1GBylFjQ7RqcRA4H66E
Kw0RctdfxYwi3ElwuUpha/8tAxQx3dz00ZKT2HSjSfn0F1asRG/PMO5/6bdLq0cf
ETfmpFL71FRu9IPd0G/iDhSmtLYLmZ1PTAOvXPrScV9BrU72X7YP7tiU6NQCRclz
LCy64Xaax9ozAmI07aX6seBiGdJtOhFyV4ThdGC79xoI54xK95zWYs9nz0HL6Wzi
w52CbRMNWFDyCCn+qn0j3R0ohmt/p3njQbeLGVtGQv72lhtEXzVHiko3fTIHso3D
7b9OTo15zOIAiKyCju1QCsdT4MqxvSILTtJ3I34yrDiwNTzRIIr61IgduGkNbI05
nO41EkWwr9I3o5Wf47wtUoAktN03bAjM9n9Av9c0SXJSHcqe98TqSAaCnw6KulUC
qP+5HL5yCz383sallKGA0fTKb2a6oi0G8nFhP6+8dd/nN/KfKYMMxhVR6bBzJtEE
akZKElk3Knm/G+ucR2J3fFY5dztaYNHZqKbcenXLEm/zwHDpYnoqjIM0XU1GzDTf
JV2iv2AHY4QROzxwiC309q0uEYfFcK8cgVtsytQu1N8/oa94FNQKzru6grt5AtuF
s6/R7pwimu8bMcAh73P53sfkuYt7DWjxef9bTlNmAImOh8yOnxccGVMCAtI04Ihw
Wd72UtGK80qOc+hewFu4Dynanht6phTTzk7+15IAR8lNi6lVB0MGAr5yfYT+InLs
gnBDSVgmUdN8Dlb2zjsK11WmP0FlyeDUr2tXZh3qVP7KxMCgl1bEJEUpfGrMeOzL
Y+/+LL/IYtDBmBtBqmBQcOr9Cp9cPoNrmn3giNtOPEQ1DbPX653LEEXHn32RXsmt
IRYMGMOhEZT2I2BpGXrwjHEwE5IEO2IgRo35dB8vJdFXVu9O5XJSX9EdTkskEgpY
NT1zVjWvn7ctHWa7g0n6yyEcP+qOmYkkNnkEUgJ88P/X/Rw3gjJaW2d2afDlsTey
oxnoctGu/vD/olM3rFx9BhgPzLjQo15e2ItKxV06jqqTftPTX/kFgIfW6UL3BP4v
7Kk8PtvcspcsoCtRFNyiJ0GtDVbQVo/fAHOKpeUCaC+cstm+fTioTWXW8bI1Qm5G
8ZDsfLtmDZ4IQRIjmwBwedpnyZs6OWAvEYEfMOVtt/K1YRR35HuFSuqSjqNwTiMc
wineEAAZQSXZfYfpPL8NPFd++TnpL1ypF+b8k+NGV2xi3vup2vagIhGNvchuiJaa
J7X8dmiTmAx/3IzOEfuef48ufZEYMYJSI2qwH+3chwONbvYldkELZehv/or5sxuf
MfiOFCvl759wnvH17B9JjP8rgCxvY1tLJPRbA699zoX/j6KvaD33Tuo6iadKjY9l
7KYFl6O4zJtMkjKYVr85MImEqz0IcHVozaET64t7mhpXPrM7cv5wkN51NPrZqKUy
/GA4hk4inqDD3XGL89mPuxEi1Ctj7OD2sro8CbAPFISJJawMCgPBToaRzmatyUOD
SZaxjiUd2214SUIbODn9zwhrLsk8WPpYIHPwrE9mo6aDafZ98fpMWQEjWsSlqrpP
AIcPUqWYsO9JntxhrWzXTucTMeU0hWn5KPfXjJarXRimrLNaXN9udmOfeDOCjM8t
49D+qjfd6MRQTWNcPNA7RIgaZ7HjgMja2ZWbI0ugqXco8IWMKJ5cipb7xevO30ju
pJRbNE+DF5g2XNCMw2bUxKoki+ttoOEUYvW5PkCHQld9X2Eq786QwU4CSb852x4T
vhugwVDDu1cqwvI2lXs6ic2ZKzEiXp+GxKSFezA8XsoxBzBre6atRJ9eK/qiYG5S
MIygcZsWZj1m15Q7qgXibZbHab2SvWizS9zW7Yyk84J1onzq7dHb+uulOzJsqSz8
dk1CYHyIwOSiD2pS8o3vnEbQ5KEh26qdG7SXuvETbgqS8cx5ZxoHSPQ+ho0/6a3B
ksnOfsZALc03cbYCu5KPv/WHuCADkdudUISFoNhM3dYHhUAmiOi+2cBrSf2nCM0s
CcmjffbbVluaIHUYvV3w2YPXatTog2OSbMq/0xln6ni6s8+6D8f/lTpmxtr8/E1L
/WN5K9WorQUA2xot7veeXALbpsWTWdDKju2xPaYkcLRII0sXXGvw17Il22V1i0Pb
/69+7d2g3QoHAbYDEpwG1EvvfEAIc40C3KDCFtVcoYyUcOm/+fO2kOx9Xujkg+fX
j7hN+iJnqBCher1Do0ydv8KslFb+VOcFrfIalDMWXzTn/4ET+yOiYsttX3qmjb2g
/lLsKDnP2McW+rL2l5JMyA3Goqy73TkdcsQD/915Q9voHQakeLe+9UTb15I0BnV0
CTsxHex6S60waqcTRgx67lEQYOxsKfwohVeNm17NvoR8LlggZwDTjEmvnSnSaPTP
i8lJ4TKghpGl66fp+Mfq57gl8gCUZufxTDsp1x6d0w4w7mO18X2TE5eseQdnoNFG
0nVnv6B3GnEkg7eoyTsI4puDej0HcM4y5IuSkwARinZBacLifR5xdJnq3gKn5k4y
+BYhPsoyYizxGj30/tAXTwyVnlMtzp0WpKRXJSkinqN0uZEOy4y+pUBhUsrETQHq
VudTUf8y9bQRcBMjcA/eSegqaiGkkQjUOiKoo6PiIsS4giuOk7YnW8jonfbLcYXR
cOt1d8G0VIi3hJYDrCm1XM6I5HWu587de6F5lBykO/4fbEaa1BBcxwZI0DR/3Suw
GjFWDuciTdMtvhSuh3fNfu+UBFLrneEb86MI1lZoaJkUbxnPXftXTUhO8uvvNUcW
1DOn7qFZtnvx3YJjXWByn1ceLj6jM+RtcuyDIDpdq58F/agHbfAQwz2OfbPv9ZmE
HZjKi9LPiEtJu364RX1xXaLsEEkUrHGvORMvQ4Q+VD4TG5gsB7fOF9eKtZ7nTmA7
FoFudT4BqhafpXlvfjmqvsjbAIVR7tzynGnTdct83AKI9hDq/xgoV0UBlfuFzSjK
I3iFOCa4QmqqJyNwDlhB/9QZUzA3+L5rCV8E+C2SDGNMSJHSC7kZssZZMxsahyLl
6d8ny5HnKYS9nCnbeKR9Vla07tKRyCpVQw1GMoaMQLyLkHmWTDB4CJh7F5ad+ZZc
8wc9lN0jD7qw6p1uAuvlAwXHwmmO8NrazRdQGR+iLFMOk/6939HBNy+Sqw81ry+H
jZUd0/CSRGSuJYpyoFVqCw1kiyRQS2uishLpTRZtAUGBu7VJIuDXBY7ncr+HwZNC
eHnNLdM4XQ+ReZQ17FdKWxCQP0JKNepdDtuLi1j2gtgLFJSjEZaauq8Dd427XKC8
8n31rolh05T0wDXfPK3R9JGwZKTSm0FzlwRVPdvd+EkwTzqIVgCLVCk+j5eMEzs9
E3yLkzpB5/nnajB/RmQkwdLjpyWFOi6uWesXcxXhvcYlGfEKLKrEVnv5oTM8a5oX
zBnb4eGWipFWGxW9DhKu0gD5qzMajcJlGRMGECdbWGEJVfToanEufytlI5tJU6la
8kMfdjhQXkIfEWv13s11mO1Xmg98wqyk/1swWOeiftGyHk+l/OYGh+2vl7DvnrHI
XU4tVDdA9YJrM0SwSK11bcPE7Kwv9NeDxqMI8gQELGeOWUa+hr4WQIw/BiAzkARt
E1fndcyYgJ0q3l3WpOHkVuoKqRMtkyLCYKq4bf1Y97J4eBZoO6DOS1ZRKqJ25W1R
hZ3ijFqOt2a7xk9usiAGWsn36Op/Lu0f2aTNXkrpSZ3lxSfNk0JV73choRUMaYvR
y7UU/aFueeQwSgz9I102k/xQ/NRPu5V3ylDzLBJlxCRxuhgkIUuoK/7oZfugZV1S
L+wKKvZrdWWjaNc3QUpYjPBwYEaDnpgfw4Dx01RERM7O7k52Mb279nt3UkyizutB
PjxrroPtehL2WDbR7B3tcu3Evn78l3MLyev5q/OmGsWoZd5FGoJF6tfNQqYDEWMk
OhBRSFsEnXNoW0O+0r8r97OMJOUNdajfwmk1WwlTB30tlGhS6/B3+UFbSwSKNwAL
coRpc+I9S3Z2Xtb5ksFMVhLSyVYPwvFtJUZQXar5icYxCCXT3J0ABwlps30Wrtom
fIqa1qorQ3EaS2Dfxod+pDRLwIlV+c41fU77jzdC9OD1SBAfJWfAurdM5igWrGcj
SKJLgW7ANksUmsOGcbN/OHlK1M1OmN23oGTzrPzliLuh9VkLiwgtt/hEAFr62y5V
ylr/N0CQsjKarI+StcTEeiF6mToxo17zaEtVP7yKKkFiLdBChUdwFt4uufpn0obg
ae9xN4qt734MS4tys1qQOYeTCUlULisPBCIbv3cmsfVlYHZHU0+CkFaJ53Sx2cVR
mXN3U5z5sLefqWTn6Kux6kblNIkRh9TBdSIFlADt0jeNORyZnnl9vyC/bQsJb9E9
yO5dWO1oV4eklb/HzYr2SV/jlqDsacyROjvXPWhYGIVxQOyF3Y0C++x5h84/MSOP
lnPlmJL+cA0S1h+YJFTQ/rck9GB57oxgx5/48RPh+0lLl9Fn5FOOTA6kZc9X418G
tR5qqX67wFcVFpm20kB6nzlVEU2Pc71YC9hxhmKATpK9wf4z6eQND6zGddFJlTJU
7TxVUc/WhVQ5scm45cUQkdQeP3s9I7hY0ARF5ZKP/EUKh8yMyGM4rPyDdQ9ld1zO
ZLTbuOQglDJJQQdtjeh6TY8dtv1yUxDrnYZxvCTIRzvtajnwiYKBBQrPYN/z6HQn
Oazm6ZZ4OvYcmuWa/Mc1MdolwzGrBse422agywxEx5VGGfwgJp9PCguA51zvmmti
YBW8x8iqrSMy2Vp/jiKdhctBQEPpwzpOg7fuTAqYWcQDRIC0itK5D0ZeOSxyNWUH
cyReTPJhS6Ndl4E7TIlqleJfnBI9jiZPgYWsxS2/6wWFiGYLSHhN90O6uOXx/YRe
JzpAwb2CLNas5FoMw3P85A7W4GR8R/in1HJYyLWsi84aMlHuYA2SlRqnbWrl1htl
6065K16voUCG4JiZ4mqcdXOvsC7wLcWgCebnJy366R1J8+xQkgFml99D5sMiLgxa
9huOwtQwyp4njG2cp3d99RWXxJT2i1CMTDHCVk7ZeZzkWnZss1BjFIxj8vnRnSaj
bHZTQcQ3LMVWBvJ2ZAfOSw71iE8M92ICpD1D2rg8VA1sgznAE7kHqqtyDiIXXTcp
yGsDFyhK6pjQ77OAOX48CSSK9JRyF4GLUsA/ww5MMCoE5+HyAD2YWV2UvrbivgYP
E8e2CMMZTMe1nT5Nau/qHxT7O2CUvMCidoBhC14noaNrekN/T4TEDmXDwkZOH9H9
HfQt8BXWVIz0llk/5Pd9CoKRDX6BrtLz7erySHmwN50aq5uiXGN61D2g5nVUKTgT
Vj32PzXT9DXWYm5dav3USe1g/LSACdh3xOmXOn/8xqNkoYOvSjDQjgZ+LK0lDzlx
oCr2PZE90aQfzIHd+ovrwaiAkdjZYGOERiMfPN0oZGN0kK6SLXWhhE0O+JH5M/gY
M1j3fSCFyRKqk38ffwpgdL3OegfELSRBupJuhIDybTSc5QunBqRvIeLOjSen7+ua
jzpUqn5iHd0qXGxKfJpKvqQn8nng32kshnD/ObC0M3RUPheYfmWle+OORclDs/Vg
Da86Bo9KYSe4PIjjkFl8WXqKOR6EnjsfyR3LO8t/a3R35Z+9MFeLR6dwYFZitnk4
QA5U8YXctLeqJ98gHp8t/su2SiML14kXlGZ66nmWs77klnNOPpcJqTEnJPimU4mY
44kjap2wDmBfeFlf4pevdTF3PIrZcFGM70S/TNnzg5ug9toUztW+c3UGYqPKn1FI
A3CXfZu7GBnz3FbjIHMeu3qq1ooxx9eEpnsNJCKA/EALwTXLTjtcDCfFhUm+LN23
3SCN/qaXrykPwBgJwnefub8/u/kdHqcT2Q2JwuYQ99Ya2nOam8/7EYf0xIxv0SA+
cfrieMUdt1bxzgHACLbJM6uHxXGrkYH1VaYoWPQI8r0NzU3FPaIxcUcmy5XmJVya
LiVRBowbBt/Sf7h4+jv0p2ZJWxfEqeOdAup1z6UZ5C8lfaukpQvlsfbx9W1wBDeJ
tJtn+wBaLZO1T189FH6gtG/usyn2RB5QOUi/du8AW6QwwVgXsBZQatACu7mqQPjB
wik5z63fF0q9XEF9esYBWcoBUutlJ4Aed9QICAuN0Kl5SgtV8Evw75hhLgntQaHC
R48/8I5qdVIsesONwffUZLRjMlZ4E2kH2WOtSfmeSGNPfhLf5vI8Zc8mQoehS1OT
s2Uo8AIBhViiLl9WNlsuoVSbF/lKnLknO5zMILTuUs3nQsFHTFKk+cPNt32vPHPf
8mQ8UYOBHqX7O+0M4ARx1XFTDNgXKkbVd/CDtd66kIc8+wgy58wrDRbp1I6CApSV
RlaSDua929l33crZJN9DME37YrRFhBKk3zD4wVKdSAygkIA7hGXzEXb7bDmG7uHD
Z7Wo+Si0rFcJbUmzyrgb8TDktxGf+zerLZeA4VxcJze6kVvnuwdMKkhA441qg2Wy
z9aVCDHZigK9RYsGSgLCWEnXSjtO7rB5tHIvwdT6xDdBYmHU4JXepg/TW0ktE23a
xXjvwzGowkrvL7wWxpUrlTHer02paz3tKv6zPYGT30h/dtzs7JXwlQ2SbzuFty8C
zbuCdsbONxKECxe9zN7ll/8jmacNXNtmR4jdtDBLqdMnWbMMRAPwwYW8cx0JoiOI
TRHEoFYzzONsi/pWcRXj0H7AfxKkGL8jL3BbCYxultpjNkqQjk4nfZJP3SCSsnqO
+Qr3PyWmuhDNGWoQIcqb7IigWfwSxLU9SPRv8m34kgC08FRCvro8/OfAnLnmBYy3
GsYa4mEyWjOtUEdgm/1lAuTzvNWAvV1vo2aanfU6p3dJiVg6Mbrfi2MQjElbUI3j
dXMmCSSVwODcwh1coyQrxNgsLiEzU9BZSi686xB0kUdZCLleU1gM83VYAgstgpfp
1JQYWE+Zc/c0S95slt5HMBS5ETkhpqPjBV9Ac/vrM3jciehkF7ZJ7XvlkRBSV4pi
7kvZAXyVlND7VODS6yd2/rhVaN7uVBEV4j9VuAvkP7dCzk5UElljbHEsmmsRu66p
U0Fv7XyfGGuAaJqOm24V2+/+9tn2Fn9e1lv3LQ35G56BUxkNNjcmoRMqQnxwgFVA
7gJmr81hxer9IeH77eLyywYhc4dI7EMqx5MPF3QoDvgTfpm3HGlxNf5bFh+/2/CQ
2l4+ZCWwRretbxyipC+Smwx9OjEVqoq0wCtanMeqoGt2EcWEglEpznuaAAMBEpD/
GXu40o7qRl5GGyoDbWbGbVgO43+yF/XX7MBmITrYi0EwmfGFSBBhUYAXDyDylMIw
QLlr5UC6mROY/KVYcIT7FNarWoR1bzQbhRFBPmE7ua65s8eLb39kt14eiwdpXNL9
Qf8xB34xAyWb9mcwTvs7GNgMSO+ADtN0vO9NXJ1ItBu0al8f/CAeYoXa/yqQipDy
OsIywQx+boCYUnSOFXu3TOCRIQEY6mHwCFSOwpDAp1TNvt6uow88K27lI7QrZ0+C
12Y9HLCVF+CkVfjJw8Cr8Fo8YBOmNOH1fxzNsfog57g0HfHXsRPRLd7Vx1MjMcu7
U3NcynD/7QzpMrVO8MOWdZojf7lKVllI+tbi5ObmYZGUGqFTBhpS3kiUE3hq60jB
e8OHwfKCMLIDLHbUtE3RfYPjChwHbIVieiGhE+ifXQr4BqlQD0BnzH9KgKeMqMkA
61bdoTpiUE+RvM2T8nhJv/bfTo1GQUl2jL517bN8pJy5GHC1/SRWyZHkb4Tpgfb8
pJ8RWHS/NpuKzcUSvoL2GhIh7vWZlAgPrZ+5/d0qfg41eHaHRT9NJZW6bAMf6mpU
02Yu0ic2AQK7sMsBhj0IrilreAGyOK5j98rOQPDgDqJPwbPPVp8VYPYon8StGWfj
3cUm4ZHwOCqM8wR4Vo7+wjTgJCY/FrOsLrGaFKKehV829AbOMtw547oExy8gEnLi
Hd4BGSCbnTJcn4IcRfLfDQaBN7YfARvV02u4Ykb2P/X7X9aA6TOExRE+559oF81V
O1kyt7YpSAS6g20KvxFwoL2dS+0sSA48HXXj0X475NQy1gwxaqsRMcLug43PMzN3
4Qxy8adtRo8onb9/pCAs4GwjkjSeVdPIuDnOIV/qSLRqONYsJswhiBCvfI1Z0vIc
RbTPxCg3ihQknId8zVByFp8WJ86wo4njQWUAC6gnKmdKg8n+rU3HROIfkkI0dZlX
o81fOJvFRC+64PWzq4r+eKQ0C4xGK0IiQKH60d9dygvfCb7h5u0ASifXeqW+wIkR
j7sH0+5xDLzaoZysvWJqjTjyQzONf+txqSNI8clFfBmY8JHwu1JZoNd7FPHBnSVp
QftISlpdH1zrxhoavxKnRXU1Z6kTly5dzNioUjGTxzyrv5UPFitVBPS6F8ZK4Z9v
+pXdvuQukwcC3NsFJBXDL6djC+ypvhAf1YCpQ+d355IVLRfhY0WW17VWTd7XT3DB
4vU9s9WVQ/vkw2Snr1BZbkMo7YigHcIhsN6JXuK0thlU0fDJPbEN5IeQx+1ZaqJr
EMXmCS3XrXa1q8SywXbeFodmO8camC1kvXR0EsDhiNa/RWMR1vc3IMhPM1Fe1I4Q
ZF7fOQELioI+8AvgFw1wGdeyJvSHZHT5HZW86iIFklYbUjcUAMB7DtEhx6ML+a9j
ORU6uFd5f9pGAxDb9WhCMoghJqoKinee0U2rbrvD6n0RXjpuk5sEWadMjGhI9I5g
fjHP32PaNIgQQ7g66kei4hodpv6SxBFvjiAXvUoGJcCeKwOlFYlR4XwcmbfzRjPl
Cg6M54RxzmNeUv9nzKbqEn/Txz7C7SWjd+XoX7Rsx+EfmU/TQdcBI5Gjv92iD2wA
5+zJ+nFNWvF0S5nMiEsGf9iIPgx7UcYSsA4GzvzjcAzgTIol6xnfXlno9YSSufB4
3Iy2RAVSNHuwzOhbazgbnYBvtb3LjjqzoWFU4QhUm+0ghDKmabIsVpdWN416qCz/
th/eYcgQUNUouNL5Oqt+9Hi2uIf4ZoO6nSaunHdLfYOlxDvZ3lSDnHUQN5tIbnVU
ptRBrBsFDDwF0n79jjdjwC/wIOkyLFQD7IgXjFYDDCZJw+T1+VZDzSrkQ0YJZ7Hl
EOWQDqIp0B99/h3njqtJITZE3rOUoNBPv/cIMun5vc/+u82dWUev7h9GfmMJfN/M
72nb/Qq9T8wQbHU32D1WpEEvzYch9Wlo5q7806dFUnYyk5DgNrdFkMkrPMhmkBj6
lHuAS5Yt8K8CmjeFMlFZEiSqK2t8M9+OPBk6fCstzB36eXNNs8m6QiPRgDgHEWdQ
pLvv2UHHWhsdO1N8+MzDONKyAvHmD9dGHdyhwy356p9pmRTnkPsbXAQIHPEsI2+7
zTfgXM0pnlLGxRYTNsnxuWoEseCLaqmK/Evr5D1x4hH6BTxWKNhwLq1dql4/ibks
dMklZTP5O900XaPAFRhmOvGJJ6BWctHQOxJLUjaeFL/4I96ly2MFsNfoWGOD15L6
E5EvB8F8jc7Eh+4m5qBfd7AUkfqfyetUlNI00WObchm5w9y2Fr+sG9OlIh9bL3EL
Z5wnBbvizkLrwGAZKRfNQUduOlXTeZnj4VRc5G3J0VAbAu/oSp/IZkuzup6YM9PM
iKPIk9+zxe+vvgeuq3kvughRBTGTduCvvHnd8V5syL+28HsFTF1rA7rjXjNoxL7t
lFCjKAwYTpQ8+dyYPAN3fK50bqkE4+7bSidk9QBnDPmTuO+iRDPXY8AiuLXABVgL
yEe7NTDgXrhgiS9YhuM7TD6ghOn7TlkV33gJwHqhSOQUakTPDujgSP+WcRNXWvlK
wRv3bpxi2OcQGG2O6iowJDgTOJwWbCyJEFHAtnyv3fw1CtGtmAVTp7t1+BBklygw
n1ZJzIvGl12NpDrDL0W7660B9awDRAavu/fLDJFNaQlDbhLT76dYxUhCNCGbzFn1
sfQ54fmov+1j6fI3Z6yTNyOltmjIYXFPGlKLErk5nCIgqNDVR8sOMgoanZ9p7uDZ
FK4ekgLp2sgmT3IdLQcqTmdSWFlhamVq1KJBPzOoaMM+0IdnE+rhHcppcm5Oih+B
qJ6DbaP1AKyKJ3T0wqLRODpL/ALRGjP1/0FK4jGSG6HJL1sGTIiJdlRuXVJuSrmJ
1qSu5s2ryN4qVynQ4gZtO4q3NhZRlR06zEuCnC+NFY3aLHqFVld89f4jMM0p8Z0p
z+sNnCgnWbRmpfUWbvFawrYA49VHKRwyl3uWF3j+aTl0lRBsmdE6+4oFVUgYIc9a
Bnxj4mHr2BqDJ0hkMscu9YE4QJHPKMAR/GigbtvT+DewiuJt/mf+jVVNrG0eYrHp
QkOK+YvlRKIT5TSJ6QxO20dwJFbYTzJEfbZNr9TZeYWoNV66OMFQoY7E/k0DkgOq
/sip2Z9M/cq1PaiKgQpf9AGunE1cBPtC1lQ6j+BuNf1h25PYfU8md4UJu9vymM0o
lZy/HXhT7m05q4aCaDvPDFvl92VL9Z2bzqZaYJgzL00aD1ZFn5GT15pGpM6hf+85
nwBC4CN+WYqKCFh6lOKx/ktg47Aq0Px4lMdQvmRU/Dg37C5Lkrxdb6X6+N1Nbhu0
EyzCuD6Yw1dTG2QvWvzPDf+2nde0jabHvVytpndYoWz3r6EzJ9EHOvtbcgUYVizA
mrsDYm1Sd6YNgqVVJE2xS5wVazVUgN7jhG8dQ+kFXhKCCfW6G3BDJsLzLVH+DgnU
JRXjsUFSPWJaFeOZZYY6OPEe3R0Neh/x94abc8AOSX3RKhvbaRQ/gWf+o++Jn2km
dU+8AftVaj4H+jZy2CDM1dRQjLs54WtXlttc5pKitg7O6ldfbqYBa5AYLM4Iw8uU
90e93+ziYNtIKS2VfGmYbj3OCmuVOzv/ZZqLZPD98M64bsBAJ2OQZFVtnqLekLFG
oHMa5LMjxLA52y4BLoMrikFrnf24DN+H6qzT7dWRV5mGo+3lcPoLnm5gcTw5O6eQ
vXbeFZTEBlLag4hdZFyHSPuXeGcCgAeXQdNxkVwDyNQQS9jJFvYG1rENCV5620N2
vlHNZLL7fYvm7ys3VHkLyyIF2qllAwIljWITupt+nmT7p9UvRiOV4oOL4fXK5hhz
r7vEawTI7Nk7c1Dqljs3Gh3S1T4VKcnWmvu2rpHRuDtepdcFew2OXcbXijtEsWRw
qJ+tyfLfKNq1N1uCqmWIuwAM6P4V+zsRFd1s4BgkfXBc30L4gaWtmsWlbAKTSRln
bP/XPxB/u6gdbd+sTfDkpibpYD1yezE2zoJytNdJZm9VSTzZ3vp6vwKideIRDTzc
UxcQtJA09VJhzcy7jkBoql9cehKGPDMCPDMhktAz9+66k01bQNxi31yuzfItPXbV
sQR1gbmRmAuTaOA2X2TJALxBli7DJl2jjaALfm7Py69D1DLZ4cYHcU5L7jUrHc/C
8VNMtPG/TYEQI5jVfol9VFPi7nE0i3p/v7RF75ZD6X4b6TzekVtRgVoX9rP80ed4
WFZuJUiosEFKz9HkPAqAFi7o1LphivuO4kJYWzgSn3ivZm7hwn6uJKOsL+LxjBzo
qWDoyVyesA5TAM/ZzO69H7X8q9nTS51g5wCzBFvTjsifh2Tp+/+05hBQdYvSvL/2
Bk/dbOOz6G+cXb8PqNaZWxJsw+b5gXWsGsAd4peoMu9H3jMWGE1xUOHGd5cFQ75n
Kh3KMarYLTBE3ibFetYicZwzq53zr6v+leheazeMDx7E3wjAiFtpV14LmCcqRqVI
sVX9lEuEuYGsebI/+NLmPSHZt3517ieNb12GRsJ8FUuyJrn/DIbkPQ5wM6Y/ecxS
EhJIFDbTYolEd/mODVvBCRS0ZIu33wfK8iImA3w7vJ8FhnKboAuxd4/DKHWHbSNC
oQ0wA+H1WUUGkF3iYJHHLOTD92W/qz5Ztms14WRU3/jjTvFlHmn5TE9q2FefirMY
ezUORg0JxWmzsQqR+M7aLBT6MA/6NjrafSZ07EcLxxKxZJMsIdla73ulx7DvvBxG
FF3XvK+6qmEFcBdTsrM+d1O0IS3I5esJu2NLFC4px3zyRcxH7vsphQQiWs16EzIO
0XAOHsAd6sWUavOjQakhmy7pWbStJvjCx8fI4AiZdbEzBuXsbCgi35Y2snhBJsCp
yWwAM8/jF2GrFLMuYB8jJBadZgCujnYt4vClLvTfIbSuhz9YYyOBBr5eRzUDR1M9
iPR138rfNBk8BqYfiTyU9wlpjO0zq1CkF+GiQgS7Y6fanjcI4f9JXoKu+LyekwuT
Ufc4qzuWe/ar+rqD7lpofBBj22p4TlhFEEMc6JsRNTWepglazu0D/OpiPv+I2KYO
7Y/MWHK792/wNxKJ44V18RKT5tKoYnypaC4Yvk/4adxJ7YblDKsXPafbOXXpAA8w
puk7KysnZKGAwjWzJZAsOfsQYklUDFiUnMhOkhJPGo0q7RxLo9BEz7PeXho6Jfpl
P5DZFR0/zyqB+hq8u2+1bO0tXoTUYRSsOok5438z/cI4ZkqGbbrxXOTS4A+LSuto
w+e8VlcC4KCr1Zh5W6OvHdTM/06q6dXZDXZVqlhxXPxYDtXuwElOMgl4/FEklIjI
X9U21JAcIEsMHfJQRX4iY6WQX2cx69JxClSMOmxlws2YcKNd/K9/Vjuec6AF+H9F
EjNnQNLY44Q1QCllP5df5xMrlZYkIeS/JJu0XcIVvJsl/2XvTtrBrtwE5FWYPPOC
/gckQfWj64TIZTwMdb0EsErbGZkuDWCYK/w3WRg+mGmjFRCP7M4IDJZHg61SBmoC
O3C/Mhae2E7e4XUApH+IWrBEqn5MA/sANWOLgow34G4M0z4UuvwtqQGY31PF5yi/
mYwK/NEhjiGMfVpLVJ5tJMbKeqrNEoDKHCguH7hNQeVCuA9hVziLmE97ImYC45/l
uMkVaf0ZiMP4ewAeQ3eCvt49QJZKUKvz5a0OAaJPVC8nXH37d++SGHYMQv6Jt0iR
C9F994eALo/lyD55o/rTVGlaBRTT2VIelKf0WiLHmMCSd1IknyxNAuySFjeecHNS
uTSbPngMMIr+rzuU0Ap4BVmvUy623BakFcQ4dL57L82muc+CcNROOdVmjqbVh+MU
WLHC/TRmgG44ioJZYmuZOW5ApguJxjibzw0iQGAnqmiztpDPwb+/BGxGPHtthE+e
dWLW5oVZqaGSVA3C7/1svGXhNgJsZuVfUTL4Lq8oTJAcByk5c3M3Mh6vS84ab8pz
piL9mnJP1zERrkFoEE7xb7i4MP5OThdxlvrU+Jhz1astLxEmQAtlGmKMUyPIv93n
tgnN5Q8UC8/NOrUczETA4/OtrVf3s+nIFqu+KNyRwth+FCIUF1xkhrftnNO3bsAT
/k4bRzu8OZ8AT8iTkcxsAOByGriqEZKYgnyvhPWqP3owlWpPhb0fe/DMkF8j82/g
ZnmtmgaXTriKOLw1pHjZJsStR+B/XFi8PtoQx0KEgDbrT8cZ/GKyovZzQuiybb2Z
WgYUzpmdXGHAtft+SQYG/GLWQw8ndPU6XmJdW4BC/pmf+lMWHZqe2xNUt7mUhxTW
sDsm0jUU3Ez9hmb99XJu0H3qvVMEeQyxIns0MGNQqKskKQLSXde9xV6E4o0jYPf5
s3u9HtnUrvyxBhTpk66y7QoWMUAcBNqyB4867/Ak0MiOyHfPumfzTqFjFp1oplCF
AokfuF3KkZZqQWEYrU59+m1ivkvH6bsUpZGR5QdI84YLV2z5R3AH6vrcXpn2nO/+
EBhtXLqCT6CUZy72NVxncPU9xwA8iEqXm0ZoA7IShfDESexpPqRog4XbI1qGa0fG
Jbd56pfqwbrcUEQmhQS/b54pRHDtgGXk7owjWq8XYw/lnO00hdu7MozU6msiwgFB
YfoSRXaCiDA7JahnJ8UTzKnQxto/z/0xIDK2OuI/hlDgM5yY2LPEO/HY0GhLPLc3
GAT/iL2bQkV2/7EZ8NAnNeLikVuI3md22eWp5W7MdFK674UM/ySom0rRPQdOYAN2
SiMOaeSoWd/i9pD6jedtvtDun3MKkfNx77dLNw5L8v5NGOQiz0flHzLX6YNkNI2l
gcH2SbE9lAhaFwbF5HDhWhBQucgADm5qtrrjzpBpjlb7ESUQCxkXwS9dFaBv9/cc
FZnOYOa0q8I1wTzlJ1RXwEN4jdmjw4ht5lX5rwPF9dwGdDSBBFOH38YKvq4pyuyA
D5ceKXhdGWAZ3wYFEWTe8Y74xHJCaBi8jm2EdnmqeP1EXcrwF2TApr7uPtyuBIV1
/Jp8e4sN1S8U3MBuGfTD2QXQEeWpbIARextpyeae7pvMdhbu6TkXa+ae9OntMmeh
nGVv/PBiImWG9JFRwVg61Dz7IrRU6L2IAMwYr+d2YzvEC8PSxtsgKc8XdBYB7geP
68PCuO6CWsdcz0FbhD21ju+raPWi/XXdPxH1TLfmCRvokaTD606YjMLrKDBxGEgr
YtYT6AsuBLdmm8XYDtvR6fmG7xq/xVNyMOofu2D2GVCR1zfB3hMYeHgG8rPC0wm1
U2Ql7bIBp7VAGBE0grkzgLY3w3s0KnHELhQYRP4P9go6yalodlseYwAnQHkVd8Sn
uiqxS83Jrs0Uob5k+Bp2UJVtzonOcQBPuz6EJyoSXc/tIIurY7E2q6LU/p5PD8jQ
85asg7mJquK8K91Zmj/6bnFg5XWiAMbJ01U3BMBfQuERtky39dFOg2tQegCfoI9x
ay0E5TW3PRZgUA4uU+rUDr+ITGrCll4Xy1ac15MrlQmIj/TGKvwzaQF7+NneR45U
Iep7sjtnk88noy18FQY6KBwxdO1VBhy5OS1FzTbXl/cgd2230sUH7TEaN/nJm3Xl
BRKtwePwJ60SDQbiQuw/tJectvrefRaYnGD0/ESSwt5xSdkkiuNW7As+UlhKawTt
Zh2wqAbVdcKAkFBBwPOK45NmiCIQtCOHJkdVwp2HZKvZKM8dwpVu/iwCj/4vNwwN
yFnR7qVQdj2svv1UbPLpyLVQQG2d6iMnL5PANjxkFJ03cnpqTkY3XrHraPiWwJ9e
fZzHVcPQBhaNna7f2MVTuuOC4vPkUWipnRA1VSbITmS/Y+SzVZ/4XBgDFDCL467H
2UzBgqkGhN6SouGMr7/Ek1z6P79mWlK7P84bcqMPA+BpOqBtMC1HAZ3FNbcKIgC7
kTKvSFMv429q5ZMM0q1iStfDwhJBHrSNRg1iu/Quvx2xKknEmTzAOH0Jf6FDGBee
XXQZOW/bpPpRFq+2ccTgEe+caJ71+nlf4ZzQMRi8fRF6X12l2Smd6YWUSeBMwpE2
YU/KsDCpm3bFx+qP6g8ofATWvsN/wVQVRFfRCERbNOhsjRulDJ32TdDGQBUkGH7+
38xN5zwhaTcHTQz6f2eIwkHLmUc9HaWo74ZinERrSQXaM3iXhzQiIhD3Fh7unueV
6uwDtqS4waizpy6AIl3BiEfNz8luIVTaHUC3nJbabXWDjRgnAiaDPNxgSdpiXWOe
STWvNok4O3UAQ3jNkVnPHyYOcWbOiQB/benbWZpMb5rFEN3Z2TDJBZXM2d9cKUVb
rOOo/iJ4DNUzkq1i/+FIPTDYgXAJf8/DtA+AifNawb2z1e7Fal595BTat41ja36O
aBIc6/5TL/8caqBKxsfSYqy154AcJBe6FTptR9D3GUT6apWeJJaISn9YQr+1OlVn
u8p/JRrDKaPvU7d9tHwRHi3tVN7Yb4vwWyaROf9jXIG84WFHjvYw6ddLXz8cmA7N
GuBmoxf/3KuQUnNy9/kVv0NLytYr9QLaE0lOtlAzWruRvxKHIZ6cMxlZAqPzQXIq
/eREI9dYJ2pXGaNj3E58eKbKwF4oD2DkUJshS7BsYVugda146/zreEhhm+dMTTwF
n8EGB/aY25k66Bqi7J1+kfj18Qgw7bsCSv3zrVcqM0cqGLmO/zqmXremNjuaHSoX
S2dCIBximIom2yYVfZ8hKBO2MZ5dqUByoQ4KHtROL2Q1G397+LYVsouG/2LX4rOD
Ynhh3V9+K87rwQDDiDUKUiH2TeZKoFdAK2dA78UClhIMyCn0+96W7t2JTYcGjcBM
6vA3jTHi3y3f+8MmD955Md0TCDRvHb7fZf+vaixWqXqMmSZYMzT2Ak179AJr2U2L
95/MrTLJxeAPsQa+4be4Atd8tRS5bZHWWt08ppKRMNNVLbOB5oOEqhnHPnSPTcI2
oeuzpiNzKQouZCYfjwFIG4eyaUl51CRzLb+2/zaLnhPI8xTCOfU+7WRmLEHjpuIT
3eN1SIBqjLEXU97C4szReKdbfeCOLxj5MPZkcjYz7J1bwD5HH0mEeQawTJ8AE3Fs
yVL/OYwGyqZhLH3sfzLkdNCucey3Oj6B3bitJQ22MLotcvDrQKU+VTnCjUiaUekl
IwUfQal9ogJkb4DUERyLmFzni4WGjZJWBD7znUYmT9wlh2BGYwBTb+EYwO5qvh+z
qefCFC7x/77iQJGKRpxB5/Ki0MjBglb7mompeN8FVGMrJLF+LMpC5HAuAeFVT6w6
43BRhfTria8F0S8cz1UNjRhefWcfdSIG9MXUT6KUCylCkD+uZllaE+hFuQwBPTWa
mJk56xgFEAbpiTbeH6XoeC0Mkuoag0QGpHRk1HUVvke8NSfcetAh5siiccdZ/Axg
uA2qD41L4TmXqOy+z0m8xKA+yMd+zVKkHy2eBZopwrT8Lk0v15Tdx36cuHay3rrE
7uNTlZDrBFi8rMxFjF6bc8JpD2Prno+KpVZvIhuPHVkLMl4pWfhDBs5R0J1nRd3F
BCtd2hOv4MDidgkKLFx4x03O1JIl2nEHl/kHr0OYkv71mXSllZkUH15J5hVPV2Ln
1wPANNdNzC4kRlA+unNBqtundh3bvP8HxKtD0ExvgKjI1kt8k0ghKTN5DJQbKnPL
qQ2kkk0ibeaqViLStFoygW4FHzeEYjMVraQw8+oH7rPaldvyt0OUe1CgVjkCVXo2
lOhcFeM2JDOTFwZcVpzAOGKIxNfna5C8TLzzCdrcoYHNyWcKTt5SzD838WqpofkO
KmuiBzL5afi1Z4KmrTh9b/xAMtruKV8zrcJ/viSquFgHwfKscdUyWhJFYTPbZGng
/sruKVGNDfMAQdpcal26vozRsgy+bXJiYGNS+d9gQL8EXH2XgQ+GBU7Kp2cSLhMF
B+p/JvOWOFZDv6mPA5zTkkfZctVXaW2VFbWmhjwqIULV4hZt8Ncl4BXhaXfxnY0Y
P0GGh4W32VEBlWGpHgC2fDQlqSRosuyova41Bk9DdjFLB5q6LwNo+bTPJJ7WKRHn
EdXBsNvZaH4pHYiU9wZP3Bu4TYEHVmE7v/UZr1on7EQpvBwNOZ1mD4gPwt1nj9nO
eVSH6XhcSs3xoBnV8IEl9T7a5XcIns5qEdza6Xr/8bAVx5v2Wh8GT9frNFpeLSQ3
xVMHik5NORmANVemHGWEnzvFt+H6iphwpEzZkuWGGgXSEzpiQqdufx+15vXzFzXB
727lodlWPtHahfwOBkdEGItlvp0xnJacqghGNKN9vkq5PmbsLYxATERRuVrD519+
cAaOlHZY5MAY7N1gtM4GsxOtQtgq7ziUG5ol/wsYcoOdo1dpeel4trzw4pK8Y6e+
ymRcooDycChPqfI3zH953FXFR+cJNUBJI47e43lLp+iqtl+kMhXPJUM2XSQ86r0q
nOmSsS4YQ7gC3zHpFN4r5A/bUyP8XRQHSMEmh7uBRiXX3oVMr8tJ8h5fek7uqm2P
N6k/ZEbZiEDtC6GXu0/g1OhZzgQC1Ge9RmzkdLNZQhGBFJDAwOUcXSqToceqfJHa
cFgTt3wj1U3nlNWXyJR9XfhniuEQI3DlJW76mwla3h9Ngw025vzK9UdGXuGOxmei
0GBfpChjKT7jcpcUnCGN91OF52JOSBaTmVBUXXdzxUVtxkgQz/LASY/FOnqlSM1Z
fFp5/yr6PXi5XCDNH9STWQB7W7n6X2igOMHdj9dRfta2a/2GEVviZhYkYHdX7q7N
n99Vz/tBkSjbWMEDFvkrNoFjov+1Y13xe1//MM6oEOMUbToUpH/IfGjx09AFacmc
V9mJa+7r4Av+IXbiCpZHBaqHhd/5ug/k2M1cmsmtoUEFJxlAApqxycTThn/gLY/w
AKAIMfHhTuEnFaNr/Y5v0bFllfwXzIPbFd4M7KqktzATMImBJuj48EXTb5dQkWZ7
60D7WS6OH1PQLw9Rht5mJcRbOcwta8ihv2E1Agb4JotDAapWk/TvAWrjtastaX5k
aYlEacqm1ywFKJjL1HES3/wATcDQ8m2V4AOOgWXuYpQFPKUW1GP0vJ294w5p6hUr
HsZNZRpwwERfv/ZwGv7cwXyDhSxpHWHnA3BIxbhM6K86FgNqjje+QSqqVJg4nztV
0899ogG4hQpEQaXqiNbCD/5q2KO2an/QglaIaPcA8K/pSHjdt7Wc29gPaZPTMtTl
8aJA+bijx++i5npSKWn+NExtihwr6kfTjmQs42HE+P1aqx1FZlwkAa2Q4oUubfX6
81FIaO4L0Pz8FBlSRKE4sKxWzwGWrD+s/ChSS0R7Xmb66VmDOcU3smDZx3jEaGJP
t8ZAX+47/cscBkhS4xKo36nnOWsVNHL0r131kPK3ztDFWDKOHPulP5Vd0jmdCeNx
cmhLrbtiuACFAK0AaVOPO0x83w5xadGk092tBNI9td/5GHIJzmEadZmIDQMXBNLw
Hqw6ZdgQnP94S8F6otAuEJjh7qZNfr1LQmirP5PkPVZjGdHcpDRWcVY7VilEp/QM
+17WCyA1UzBGCJ/zVFq87ok9Jjxqx27SedIk+TUiQUk0Sv9bA3QcJFFG9THxU/WF
6Ck+RSDL64+6GdY0+nqV1AX7unFHufGvHeL+gL3FxvHbUc4AUlWFv8bawaJynJo+
FcGnLhazdDdRIUUN39GQKpF4+dBf4Vv98BKpXriQ6ZmKjRAuDKJzSEQjX92/HE1s
s4NFYlKfaWMPz7oQbYp8PG2+nYt7ziuTksm4A35xl6pPMDl9gjnQBXLnPNSQULEs
jOi1acrOlhrsDDhjPB70O1OYOiXf8TcxgVgetQGCXGKkHjbaLF8qb43af+teZY9+
K+6OUuirIK4Vbz7GQmQiYwx8glYYHVVdBbm7zsXLEb493RqinzfDlAbbaAkmTaiJ
yxr6MNQKV0FGSQXMNNi7FftfULLncT5oC4v2uHQRxKAd7DUBYH+coHI89AvVzi5K
sgck/xLczViLNUjzHzubEkQBDx5OyA9hr9wb/tGP7zj4Gh6RWz13t9oL1xvtYnDv
nNcIfwIBNgo9XBenMkXdWcXftxkQq7RNZSkQMChPaeFMm15YUV60Ytz7MQ+0pEv7
myJwGo6g5McryTwFm/oHnuQu4HEW+Xg2EkP8U/MLNTRO9oTDusq+Lr4HzOyCYSmC
8501kmstJ0jxormfgkpNDjMQq6xyZsRjmobyc/EW1QRA2IU44R1CiyIseA3+qszK
g1KS4f1FLbOSMQaDFrPATD/Tqx9bLie/Hd5lDzJQV+iMaXE8Zrjk3XHvU3ev2Vdw
LtiIuaM3lP3H7IFlKfr49ISYSZG4JvkFwYKkva9IQ6I/oWz/oco88nXAtqeaw0Kb
7BFrsFZU3IhgiiN+33uyIrYndng+C9qU3ire+vig+1Rjuzhe/lx5QKnC3TRRlqWg
FxBaO2QSTSWqaeuTMeY/hT/RwypCv8esBkK8WDnwmG1R3C5z+7tULy6i2JxEpRcT
If1+uciZguKRpI034GgSlIENL+ita02g3Qwzw7kQaHl30qcL8pUrGPzByJzndL3H
WtBb/5mVs1RBTxFjlWsdgUcQ92iOH2+Md0/7U9b4ZMZnwz4MikxH4y3tZzEL6ewN
K9Vuoyyytdt3awUkGTldCyelzGbf8XAREN7BV7gvp4oAUfyl/Eh7o+J34UtNYo7g
ZSMnAWKYq8Y3YF9kmEn4rnn5NaEfswXlwpWtImNYqHJtBFRp7Pr7NN/nxdF0e16z
9/mjoMK+sOElnS4sXP8eWOQ1qioEIJFsttjVXqP8WiY9m74fNhe9EJH9y/glzOfz
tdS4WYRoJ/2Bzgk+nEkBSVnnaP78RebcKi5yFUezou8TZEDN7FrQ9uzQMEhDsOCN
dLWgd/grWDAvYzxQxKEekLDX/F4oYv8mj/tHyaiha9ATB4/84OIheU3r0ai7Yxpz
QyQEeTyB3hCvJGYcnroVkkC4+dWBSzfQIvR5flHf7TWJn2hZAXHsuM5Ytz1fLTZ1
cffedKzg7hEh09ieg2LiUjQunhmU1SucXJkyCjxs8tX0WotX2ntSFA2JqR4sYczB
zwLFOS6/Qh26CImmIWlA8/XR0DrG1bXRfM1fJQTyMR0djMN38k51bKp4gMXKjPFd
AStsxRxlYKrL531mRiZT+7M2aOzgO6WiaXMQnSIGrXg9lZ3WdNhYN7Z7R984vbvV
49fUuD8ZmibOgkVoP7ebIWyEfv1YBOYXYdaxV5MF/r77T3ZNJGz5zbJqX70opXEn
tSZzgV1eEfCop/flVXRJVmfcqOyluJ9OwmeTOTMGGJOf9H1VfHBgBc6RlDKjDFi1
ZLss+y7dJJo8CWDOZuZYdfkTlXFpnL6IVT+jv7MtWsmSTCwSCnvW26WJ7YVsar2t
cL2G6bDFRWMW8wQdgYI8a1Rn6hvCbiacgpKFauXbIgN5NYJx6WLHqmRAHOtPuAKo
IqAzX9AcqJiHY8ErXaW1TZ4Pn9VWtnYdygp1+ah64QsDGvy96pOyqos6LlYXqd6t
dwVa+2qJI+AgGtD32ZokRFkAwq81QIx1SnfVKT5L2KL2DKqR1ZhIqc3Ty75CnpWb
yRqDn1W/68v3qkIVyMYET2lmjFNn/7SmRvhUR9pJulBmec1KeukGbv6KinCdccEZ
FIm4DB5rcSm6WDag6/Fi+6gh06pbXRiqOGRfkWa77TlAtsS4xzoLq2UBOy1gPsZl
wOCdP78DVI1e8ylFTazniK0pjv1tw4KdqO+vJqJF9wPFxncs1UkKztPylLGUUt4I
8f7UQYAHlLdJUX7HxwFXGKGKQkgyRcFPP5idGgzFrvacz4fyOdVPrpXsscbpGIjE
8ggvMPxhrc7nCQUqGu6aO05VZAN3gGZYOsGMOMLDonUh4bFaAPwwPAeOiS8y1FgQ
tuZXITpptu/OY7asj0oZC0bVTybW49fwfhinOpVOENJwzwz0CrT4tlP/k7qaUpjJ
1oZVsA1w4T5jvNo3FIrPQyJ+lBnyKxLmzuKfmEz222SnN8K5XWinZnSK+MpDdT18
179h/neIpxLjIhUwz4coTscP1MApBJpFkrSgKiKTasRU8OvMsGkUNanDD6iuNpTN
Rp5G8NAb08DHlIoM/Zd9Bv2ra6PN1nrJ9dU6u/FoKblKpbNOQwDexKTy/jiUBOsW
Sy5Bg+GTfxcp6OHOlIXZffYvl2ZsUVfVybI5zQJEb49A3b7szczmS8kG3sTan8NW
FAz3msZmkwb9R4KlrZzpxMg3LdtOMC6XufFY5Ut8XWznl19H7JFIHeGg0ODrcO/f
vGqUYDYJAzYq1c4aGt57lYCXgdsJaBakNQUE5ItjWL8I99w2/JyVbh0D3nM/YU9I
WJTAtuDdeUa5UKR16X2QZ439vc0sYCoLg7q985yJAsNXKG7sozy4jWTLKVmwTN8a
3ozzJMKhO418I4dLJYCmbwq9jFGw0g8CIt1cnqJ/YyWRMRugI/nWvx6PDXGlcutJ
CKpcR42WLJliXI0gpCaZTAAx2QzhIUtOA0xJkB9Q3wzqrN6gP2SqUaIZ9IFyX9mQ
KbJcojnlB2WmOiAxFQuTBLRR4oig/Ctkdid7mTlUB0B5WMAryD2IKg04x4K6gAbq
xxpYJNPOz9SjzUxJ2DLZK5LKgEaMH+ADLgz9BxrHguOGeW0KOjQIo4uK8oKLHWOJ
4TV7Ii65mEFeSNRq1wNoMtOZk2yEV/R5oUpk2yr+Wkpp0dAjb+k465YCyFUdKuon
SkbZ4e3U/yKWXibk3QLWC2x5ygWTQlP+qaV4D57hRuR8ilPLatluvcfzd0h06z6l
sW4NsE1x2DJ+WRyAK31EwAqq3vy1oZf7bopYklfz+PTOLVsmxTWZvZOY1RW5PeV9
4yHHyL9FwBlBQp19FXmflzaJUmGiPNn98W30BkMQyB4pKaTXZAjhxXaj0ubrgILz
S8m+15eHHT9VfE/DrdsSpYImz4hNsZyIGEg/Xg5qZZ/08wjlN5A7qsgU+nH+k2IX
mXbgd46TqkZaRQCXlijAtJ3BBc0q+7Gmnic4wdu7wVtSF58wFthbB+pZo+BbPN7B
j6ApKAFc4LpWmnNjKPuYpixcii1Vc+WpXVkvtjQnzsOvot7Dh9F7KuLedkqI9aZ5
yEheDUv2uVeO15tFeb3TzGH0Kgra7rMCDgijaN92pLFLhxkFRagqZ3l0O21JvZIj
ArUPpVZREH9piHWdLaowvLP7pjEH0jIM9EmYLMopCOKHuiBIvnEHnQBP6O18VFrc
Gg3JdTGz88dlFsBisTlPmF+sIIkfcktpOxqWZiw38sHFexqurPdZGnZil2cY2aRs
mVBa0ke4ajD3SvhtM6Xs+iV51EOzRLO/2/4fX2WfMaFaXXCciXImZ7jeYgV1HVcb
JMJ3K7HOv37ndWIkP0nUR4r4niD0E+zNVlaDyOKHAcqD51Z+MTKTQQlk3bsdPMU+
/mEHlEa5rr2uJTxWIdJVweAT9jd51qpJKiiSiekeVAtRo9cNXaiTP37n/VPR6MxD
KaiHx2eLf5j33s/Zspp1AMa/v5xbVABmOQLsmFDjZjji8mX5FJUttpsv9/PRlTyF
21MpVsRdXcy5PdrS+MtAD89Q1p4n//Ha9wvkU8/B+uiwGWshpSSGobUZceED/jLm
ijBNr6KZE+7nL0cOAPqVaVUe4vKdAsnfmlHEB12e1Kq/SZ9YB//VHrt/msZuNLTy
A4YSolgEy6NRYoI5hM+gMXgdv38NlUj0IesozfrOCnqPF/wUqHDyTZMqCnp5iHgK
GHHq4lIBV3G689LZClZZ2r3UNXQyobx/zWnmjbDDoUOJBycQSQSWgZbdt4acnBy9
wx4gzFH0br2IPPGa3YHYQmySQKs7SoZYwoMwJBlav41Hd2Nf4nAkOpfqWbmY3AIA
JFhZKE5weymHoadPHKnYy2udBCt0zE9bYbvI7BWAIkc7YjvFMmEljyKRI6cQ+tym
u89EzpfhnrQE7JSSd5H6r8ZjMYYHp29Eq4o1/WDaG8E84HEpHOoPZOhTXINtqJ5g
I+jK2RXzfcsrGfggTj7ckd6msltTeuLW21drqDkRiRg5bSNOz5FZkd5Q2GCWQYqW
66tEYgHx06GiJaxyasyGxwK9lavo1J3N52FSZXNsvf1iEmwUwVbDuhpdmG+btsop
SO947PnWMRXtjN8Pm8AyjqqVVWMjuCWj9xnqgYe3bXeWcqzkIIHM3qh09OQn5IMq
9P9oAmWQsiHVFg5VYiN5bCqYVBg7qRxq3ttjcMcfWdXU58PAdn4v0bDFJti8rUqg
8fsVZd1CWSgxphmSrFgMQLtXuSKHpgmwXL2G+lW3vWAH+G86C41+IjaQS4QadYGA
LuSv+uDBbJRTLQbEXQloBl8lZNfzZX2Q1m/UK155OigNb0XL1U0qlfL9OqPY1ytW
hzO5TvTRaxrltiE5qen6cD04V/Okqpj1EthsJgPWEhMxt3U8fGDpEw8/P/PoPCrm
xiOFmXqX/1EA25UbGz87cUXn/nRvD8GZZBt9CbfiPGwLt0gxzbtOpzw7Jjfq/Guh
+4PHAdp47ljTJE19vqdwVmZwUEaxyzjcMO2RqPHcdR692MOiA3vuMQlzZjy/29zM
qYq1Oo9J/1ZJIT+9Y7BpQPq4oD9QRaRgwkzg21WfopEnlzJFQS+XRpooKRyr7U1g
56oz6oYGjlm1tx6hQG9tnz75Yj5yWB+vSirVFC+T+0Say3yuFkLY0nmhPO7o1Jbc
qSrLpHv4gIHGz/jYCabNn4GLface23hW/D6HenwWPoi77RNyYBPY4cOMjTZQUvPk
vy/Y0ADcXGUv4oNdV19T6mUa9isblK8FHTQlMdX8e+LCyJd8Q0+OWiJBLbJ+CtgJ
ZqQwhd7OEM5dsD5hyoIWE/lowt3XPjmofE8keUAOT/5TQ+SquqQFwuxcfUxdJAzD
aK6ZdlTXkAHlN5O8EdGVFiyxxX5EK+oElaQ7eN34tdjw8vaqyFx+bhU0nTzaTWi8
4ggnGDlu6cHkIEEpY4M41EBCEzn2xsvxloErcQPpoQTqk6T23GTXYnNuR4a/R5zu
jQXAy11LE+8O+kceSh04ygiIhH99KHRHAcvKXiSmNq8zl8bnru52zPV0WZNh275v
IJTul9XqtJy5BgBqDQYSvA6csBEX11MtvUMDn6s/d33expFHJgmzCbbY/HG89Val
v1aLzFkgTgZdQJWWkm/0b5J85DFyvLJBYFgax+/Xr2jJ7Gdde7drdmO9YyASTKmH
kBnQSrZ6BUBKXAlqwRCqmmmfZkRJvp0FansUdsDVCWIM+jn7hq7Tcc9/Ckavcklu
aMnxp8U/T9aNDFkZ/kYzT3oFedOYaG5Oph02u7ljUv361h92mH5DvdSU0G3dRKsi
bX7sbhOUMul9aAcQAA80etyEQY3g2f11tYNs3kRifEbBDhEwQ+inAI8oDhta9yAs
uG+IZ1yQl31+4jj6APRjNPaJMdKR6QHyYV0Na3r7J5N12+nSCrc7C2C3JV2i9qkG
fCaJ7iEvMVXXO50MoxGjKhhOH2ppJlsqIwDLZZznC78KV2AshuwMP8g6e3CwK6QA
+X08wHHbhZQeXrxPduUj5QPwOaf6pgP8NtHazK6Iq1YBykLRijA0F32JOCQSdW/m
I1gO8rKRLwlkfIXItXgFAugRQqe9FkEjKBtlE3Fyb8b/fP8FdomISxb1ntRR/rgl
icndAbz7VnOn9yl6SDsTIIxhhyRxYZXjOfzfYQMEusIaOEn+vPbHDb+pqjQI0B5S
YHgFclvpPjfrcG0vNSBM24k/HikXoP+R1QgfhhCQ4uLsh9M979Oupekz15wLpXrT
ehqpaQ2Phl/lbASFW4mUNvNQaOj+NMwf5U2Q1QPQHqkmOhE9BZDgkRkGkb84ySA1
7rXixmV/8ieknaWAk/1OAsmC4f6D2n152FKppvqDuhJx6Re46QAAhPqBWh1xi6nv
a5GBdofPhi/WBpJTV6saP4Nfenw22g8mxS8vjBLYXljrglDqvATAyc94rlKOvvOG
GZagOLbQ01SxMn8hdJ6iRvmj8G0BgKINndjJbEKV5DkAv5R3DnLB7uqX9SWLH2Y+
B8zB7LDB1cww9p/+DiUmjnC6+7j+v043y67H7DHoJN1p+9SeUAoV2Vllp0Vppxzi
C6G9mQcqzdkytPKlzuNNP6bKN4CjfnqzIKW3WLlnwNpCiac51V8Vyk65yj6KipN8
sISWf0SyT3aK6FvnOjfK3c6NxrmRrwP2l9yoK/f1KsdfTauySiuBCJcL9iVGYr2l
dTBffJX6HYdmOtqXhIFyvRGXVcGvn35q/pVrbcDXZt14TsOBFzhieGavRh/qxNJn
vj2X/u6lv9zIa0OfFjk70PZOFWQR9QmfkLQ0XKJSr3B6diWjVuiMHHusKyiGs1MD
mLSbrmYCrBTRqb/H/0ZA1fivGFv9IX8319cGvzIaf4ailNYoQZiQV5BVZxu6DoV3
Es1rcjeEl12fZyMzBlqRE3OywHWTyLB4qxwAXIuEc8VT6VD/G7wY9xdl/LZ3fbbK
HyF+KY5c3fe8E3D8dWOTuXFNHUv+agbOZ8WNLqGg7TCdiFSIY/SrvaGdNhqTTj2W
qZwPJNHZWNu34wl3GrbdmnfoO18mXy0gsSqeK2ic0Aly2wCFu0igCI1V8aT6xkcC
q0WHX107gOz3jStCUNtCB/THISyIfX73JG82vVgnuWUWVcgM29wTiUKwrc36vSz4
lf5AgGbfhOAQSmKlPoZNCrwHVra+kugf7oqzYtkFwRZCaoBU5HEPvGClHpD1elwJ
PDOvSJMXkFGYd0MW0Arn69MEcOqvLeTuTU9SPMdr8bQpnkZCGHAIaKvJImZQAiCy
9PxuxL6y+eVBRRWlm+yrPDqzMJGZXfLqmsbtOEenZ0vaMTGzu1+JQYXrncPAwdm0
hYmc411GP0UZhIRvTKPuwMCPXqRutn/Kx+D5K+rfr2tn9KaVZ5bDJE9SbhcyFXAI
oMdoOPghjN/Cj7hBZwOlxCEFa8JuzFwJmV1PPluG5xbmKSbwZ24iaFwe8KC2RRaQ
Hn7pTz8J/QVxGc9Anmn/2+EF7PqkL8wecmf5tSaLl0ECxOqQNQg5/yb+JnjiQOEh
gjqKy9VY5tqV7erM3Bea24z5FUwlvfkxXbF3H5328S35cS0wSlYn60wYtTEJkqFs
VKLwCivQWShhuwvof6e+dYuDjPBHFEOHkA1DFH/ZPGjDa8yEwiacr7cohU1Ez23K
cnVdF/TsI41dDChmOKI0ggsJV0EvAbpPglbko4ElYIzjk4oF79qR5Q29B/fps/tK
AgtgZRjV80E56A/sBRzoHX/f4gZWWcHp8OIcSPd9zK3zpfR38+XpWpg+fPtKfL8Y
nYtoJ1dqePiPydvnHCXJqAWiYAd6q7f1DDjXqugJ0yguhnFGhFU9oX1tHReAUaX5
8J0e6dUXuhcyuzBBYyGaGEgikTPBmTS646bI1Y1NBXgi3cCW8DRUOv/Tt/yKkHWz
B/mwC+4Y63JxCek3noCCR2lKw42ckAosHNwPl10Dm1ANEwBMqrvG0NWK/mRVOxPU
IAvLAFZ7Etsw6WsT0CYLrnPVOvkWN7tujx4cRCI6o2usum2EY3Tnv16yrH+aH06r
2ZioaKne6HnysC0vNCY+3l8gccfsqCT9x+mdmYbrxJF6dPmlUPHv2yvS6fq4vQXJ
0qHzN1N9wnuZDi/63qLCc23ouVDXC4x/4QtQURVYpASmjUuILgVz2mbT92FU37iu
lc1U3VfJdXnoiZjkMnHMV4MNABY2f1tRHBAYoREykA6xE4xA+gjaRJzj7BLh2p8t
2zZMf1WDikNeX29ISydEmDyo/CRDdf8FkUTZKHk79helthSp86i+mH/Md1ZksbaJ
iHUDSdlZP5Zaglq7vkS1UZ8yZAnDPoa2KIabpGkaKHNYJ3rTwsocQTq7UPCa1s/L
PKrD0ItU/Pylk0ZJu03avMwge9DgHomYH5Kr15Gn+6vO9Thx/rYlNxLih9yrt6dI
nRgcBbBcK6/IQ+iHHfCWDujvQEvr3TC+flikiYAJXSTnH0zgtpp5MaX7uV5uuR0A
KQWf/Tur3fRFNT2fGRw7UdpCArWh05ge9S8uK0mhB4JH59XuPO0krJLMEHPizP6F
s3OSl7gCgnVk1TmB81kily0NDGPswwUhDD9XrBlHtIRvnudypn7qZk9lHoDpmMMy
/pa4up123xO6yk3ruIaa/kksFp515n7WPvZ6mOxgWDQR83jamcotWL59Pc5zjnLU
VNpmrSJfvd9E40FHeFJX2wcH7gGUi/w37MSC0iAWR0W7+Vkh0nUKZ16fNtSGfpsK
yRM9tcbxrPYoDvB4vZcpMbEKXp/TmDab/OGIFQ9Twx3z8UBA+bLF0dXhAav18GQV
pZKTij2aG4MeTjcuZaOfDBalH2PPQYlVLEyrsagK/EdoCd8LiOoOn07IA+X7aX74
Z8qDSAJeMflhgOcMp3ke3mGyBVaJeJmW4uF2PUSDs2Ub1oXvPeIZaNPn9xeLcbus
ftmSHfWQeNa8IfjQMyQNOHZffRMwnZZRdt8iW/+8uMSe4mkuaP0gB+V1oHqMX3Uv
YlBQwNU2Rk1YfK0WKOnhJp/6fKtTNtHn0UoC8ttfZYyx1S7rBwlxtpqU3zlfRajs
q15B+Ca01ZgPPrgXUjsU16CdOSbqqFdBq7FwOYI54EHo/8+NiT6Zzu10inYR+WT6
27qmRxKhZwKSWbGEgJ5nUB7w41wVMH4xwI0AdbSmqixRLfP7/l8w+SO4XCkUdtbf
eRwlJ991FVEIIerhAE9fagMqaeLW6ssBR/+UoZhPCUYpIEVUNaugFU3dm8ndQpjA
NfqOfo7SC51FGu+/5CICERXcr2Cz7oYrFqUAcdnZkzBkgt1gENPm+usZrNMw/BXo
KkB4x6/hRwLlJdsh2VYDKp1efRX5SBqaOVhf9h2PGezWUhCIydZJiEWaIZd89ZMj
KeS95S7UzQ1toXMNek46cIFBcA2U70Sz+56MvUGa73UMl46j2GON9pRJBqynxUfu
huzdilUT3tBgg+AUj5lFhpN/rlUXe7zQR8tTOpd1bm3BdwMT6/K6MpaIsDYekv59
eb8UboAG9fMHBum97T4TyDrJPvhcS+WkP88o+Kf/OSxrqIpz52wcAqZMzWZmLcf4
cQjQwUNSAkimgxCMtCqCwRiDDyotzYZY2CzbQdh5vB70Zl5zuYzNPH6iwZ28CGUO
RaPtlP6l57OBDx3qzRfK2jBpAyzQz5JVuORM5+pu8cMeKqsA9AUItOVjZlzqFpXG
Y/PE6EV3rwN6Bpe12L2Aq1ai69voNXro8/XwR1VDAWpeDE11478Rm2cRwxtS03/e
S691qER4efC/heu5IkE4+XlCaZUfWvbZP7WB1LrHdhoMGZWrAApqK4nmJC0z9T69
L1EaWg8HCD/IgKZjz+oZsJ48WCqBrT7UpoLoBVQIPi9rAa/HgKMNK8hZfaM9H9qR
+2WboqezhnjgcCYaFfNnIPJmkfDeSIonZUyx7JEtH2I8GNWR6k3fqgSYyuz7+CfW
1p504e38m9ybUcvseb4ZbQk23LbpsFb1usFJtkhFoKkt6OjhRF0Awmq9J0gfMNKa
/ZdqfEzWl7DHJUwH8Tw45aCRlIm+RR5GqyHAu16vl1+LAvFvN6ks8gRobwuHDYsr
qTn3gV4SV9cZdqPk/r5YpkIvK/BfCi4whVWejix/RJHlbkKwl+/UaoDmk0zhQ4HP
6bJlIzxZDXgX6EjEwhTglz+ROA0C2hGqwps/BWuIz1BbVlKM/O/GSxv+zq/RB2c/
08rZER6b0bXb8L3lr3Zyb5pG8m6pkSwfspvrRCOlv8LQJURMBxcuDVBc2ib0DreL
5OUFDjZL2To/raIFSAYaEReX67S5S2Z1JM+k1Qn76tLQ/j3yZxBWv/5RrIiCa77H
ELDNHVDEde2hPliKm9nlq+LzkvNURl58e8n7EBmM56v810UyTOlKTg9PDg8qznoM
2Jjja6NQFJ/isLo/Lyf9+JpfRetwvScXDvxPm7OfmCfPUiGfzOf88/MylIgPd1m4
Nc9fY4zlNjL2LsE9DNoUAejawhcz/Oi5AGgZ4uH/+E1F1SfU2ERes3wOk+8lw+yu
rHhyC7XxLJrnBny1aYMA4xX+3q79vOhGNtKL2naxWlfNownCy7U6ODSt0mv77Wzi
faev+yCMXooLLaefWGiaztrnNsvdM6Abh6wT0IPpQ2s+XCgXgKmZf/GeNPCppaP6
dyzXO1QWXoTacF9vhrQQJ6NBCnmzSYWYvlawMqNi5uNQCzRp1fE3ECOQ5nRNBAPz
aEs/co/N6phXbWoj2ug/AQysTVNy6IFlI5RuLif0aYIE53PZ3fNHqTCDuci0Ahmy
7cMJ/6tDApyE9PCn5ptl42la5PZoco7Z2Mm01glGRGcI5tOhlRjd8dZeN7ENykgc
nh8QiWmZJp8PatsQNRTu8dXoO6TaPCNJvxRJITgA8f0Q/DWqO74lrU/TGPOPWfT/
FBUq18vsgsENxwmZNNN9JbuL/ATQqrQubNHtQTLEU6UrTxXfOOCy5JN0eYZjlCsx
t9Uqgqz1W3nAmuSNAN5TCmXAUrlUtbNw5pR5QHyDoUhhhMvw6c/GRd7CDKEEHGPk
z527RdujpMcholUlSMkJG68J9U+dpku1ugLAjtQ9ZyPlDFluI1/TVOmuh6jgyyjC
oLKKCgGPWuKirQAdjv9rD8clJf/zWxbMLqP+8J52xJAHieXE0C/Tp5o95aqRmLBM
xEWsqqN+WJVOnIBBNzv0xDhatXHrvIl6giMiQSu3petqZaYegjMpxLeNu+oEFh45
JyUef/eBSYLVO+VOg2DuehD+3tlfnnUg576yQjWU4Elkh4TgQw7AQ9pJMBs7UFR1
bo/6zxmQCDDnfcQmViuma6mYlNgofpHyOI76W5eoJMahhKmHxmh6Q6jkBMkZYWEK
LDeTn8a7jHUKIme7J//UwX+DyzBJDWuD1cj8ylG9P+oagpmrewov+fx35z6JKkNf
MQ7gMXBi6uFNOHfLRNKtwGVupYVL87LdX/M68OhGBS4kGKllv5lSX8XMKbdSmlr5
J+cp9bLooG9abE+bft4dP8Zxs6vDBcpMsjYQ5vTP9bgUDtd+PWGC0j1dwRlpDrPl
0NFwwi8y5uw8UJkZcRUfzqRev80grbrnKrZ8oUeSlWcBzIMwKCYDo8h4Ito1gKw9
YnxgGoWA3UyfgiyDUR0xwCtMO8ltyWME7mGrfP87HVu9hQB4T7wMVEqlLITI2rqa
/RVb3nPAO2/dG53bCoxH8qaqwsapreT8Aq+9Ypl9HWH1FqKmfll2a7jdclZZ5FWO
b/jB1Uy23BJqdVf3AvxAAEKYtWji7WY86HDRMJteubk9z6L+Eh+eZvRxbLqoR7Ut
9/Z+D3RaQHF6216pOscq5Oi0gzPqlOuH30ZoEIbzCrDtKD0jxKSgxFoUnNKe40Vt
IQUkq8LTNlJZ+haXrhKqoXfwWnqRyQNfyujv55cmKIKy8l4HgkV1nqnZ8Wib959b
KPb6AuUuZ6f8JmV4lbfPjf+T/TOZvDuUH+eHaHaOHOlXhfbvGjTdKsDHMQ1GbnDo
5woypiwDsIqqbsXXLZgPOMp5m8ojP6Zl9AAC5rmjOQaqc4kLKme9jnhNDkIF+5Ne
xQ1ZH0P78iDIaGicO66Me3R4cGXAXzSWzQ1Z3tKyiQ/OoRhUQhVgfvSZ5gQaQZ5Q
PDX3tjkXo0WdPv1MLjk9QOxFLyk/1uzT/eBgL7Iw/QqSwCZ1AjR3WYiqGsGJyRwE
FBC0q+JqGgrNdrkfPVXTT9TY9QYILrnhA8Z3Z5HEpe0zEJE94kFsEiO3n8Ilm8xz
2i/k2rUQh8HplF6JxkOx69cfeGVOCAtRy5OWJayoTHI3NWUlKxyMVTxY0TQOS/UJ
aO/YBq7rqz+39/OhHKoml+yXlRxgpwF771WDAw2V/RwyS+vbohrOGHfq1WoXLApX
lvBCp+uuUiDP+Qr4QIN1GPkkaBazf7oj2wy4HSs3mwo/fiODG9sm/buEehN2TuwU
XP223kXacn380pF+oRzyZUpPvJr5hpIiF1uD4OSC5lyxZajB1PaN4SMMjT3rJbK5
9ahM+by2XuGBPJ7HPrR2qk4KXUcW7Pgn/Ql2Y6oqwjGCBNYvDw9bAFqQeV1BNHxI
/eItXepTn0uxokRzGBxrXfKrOaIghaKamlvwR/tkpJmY4rN9QEL1uYEKITY1oaPG
nCHzXI+z/RQEUZ7y+0MnXF+fP2/5jklnGa43CA4cy/iPHpVoMjRxHueIGuBNLn+r
S4d1JIDUwRGOOFr8ejzu1/fmFLsDKJVFu/OULTVVSAgv0IyDFakQI745Tur7PMMC
rRV2tYIVWH1q0sXTEvtPiAxBWUxXUwW4FxXWi4UGcfrNOG2ufthDFXyfJP2klv2h
MStOZsYo9wkOVYafkCAYZ5T5z5ocxeVg62qYw+waXnllwlPqHFqgaYPHk8v1rG3k
VSn+crsc0EjP/fSdT30zUyH6VB9RXfGR/c3mXlQw5j4n/jYCOwrunEjauaeG9fdg
wgqtlKpgvuJQWzWzbi5rQrr2hhtX2xG4jWMSwO+5BsiAAzWDsMZycS8u77XbkMvR
IAiMmjbnL+Pacg/p4x/zJfJZb1zHYtOuEEUCbwzPYFz+VwhLJY4F9YDJrEDkBUkZ
yIGjwrSreOu/DWrX52OGyPOdhrGMj0UXdehLJqLnqtU3gLCrZsaVpTr9gks8Nk8W
etFN7mQSGf0vQ34O3dF2DIauCDD9/yPLpbCGoMCU5e+TV5Er7ocWiGrmcl2zNQOF
1YISUcShGzJT8rExdFZ+12E8yl/SjXmk191pP1YgZe2zi65j16rwpnNoVHPcEwzi
B8uBEkzP7L6SxoqrxaBEQmvJ9Mt2REb+IrAL7qH39CN+LAtHRt5i4+1pHU42eKq8
VbS9YA/+gF/K7S24bLAeG3j0xTpl2jk5wQwGhu6ZWuN+FUpUqN6bVhebXfhzAgZk
Rs9iVZd5DPHljvB5kT9J9W3isl7FsURRXT+EmM3oa/0T8q0+1IZZ1XjNu3vcfZT4
5W1t5IN9GmiZ5F9FJeogT2Js3FY1ZKz+2TjDkNH3jxwKzRfrtleQ3Fyk6WZUE3li
rWuKTYyOuVkBwqdkVm02KxL9tTIbnSGRj9sNa5LqR0Iq2Xjw1PImj53QEFis6CyN
3kutyvT4L2gS8J/WLdfQNuS/hghLb3Y1dYGqpbl73M7PXc4NWJPpvsaLuBqm3XVt
Goh2fCQ2XBofgCM2iXRUcd2mQYgK+1kWOhuBCPGvSrROvdVa6Fpow+TtdcPQI0QF
b7o18BFzXubd97tCVKfNiKs8H1yK1WLYJqrCXzzyeeFNt/feJRMhapdQ5/5V2w3r
yuBMzyJwpatdQjCmQO1h0uFQIINGqD3AJeR/eUrBjDN3p/XMzA41Jnxt996V2fiN
CcfTh99S1BUZnczRFQvOROQMnZ/9hWRAHrXBNooYMBwk3HHw+Dr+cpm287Zj8ul7
EnyewjlM3PS6SHABJ3NypHROVApdsjAYvawEfxDvN5kSRdeE4fmSCEWN1b6k9H7W
xsESFsk1xbPBMwC71W6AczoqESkHJeOwfMYSFTUFr9nTMkTrwbCB01ds7TQcmKf+
wUEyic+fjOyYu5LEmp0ZHTNMauJvyM+HW5EoL+kmq7CG0i3fVxkkgVQP90EztT4z
fLJX5z09/91co4hj9kcDz6D/5NL8QltqLBaHBXxctPu9CCu9enUTBX3dJIi2EKr/
qvfMP0dCI1agB7YJGD/NbXFfcFDuitJ6OiUlHWWXOvE3zMWqvNkuLsyw+lA+LbRg
eZps2jDlf3P3aJf8D4JrlRRm+y5JTqDavmoFZC7NHN63A3lg1VJFsoblqub6iaV+
9l+45jVkrVLNO6LPGRCogQyonda7YZ130YCUExsO5YCjruer4lttucSdO+tNV+Ub
TmA4PC+SHZjYBHX6ub69AowEQOoHU8i19jHOEn+w9qE6819MCIKbG11KZjwKr6A/
S4yuZNLkMlUc8tCQ9GZZ3Sh44W3yCRgOD4fJODDx8FWTzE6nKVIVURrYApsHiBHG
rT2Q/wIHL9dCyW8QYCnNGm/XLIkzt2isAMLQp491cClZtg3dm+JS/ptuja/B7msq
p+Kz7Xecj6bUEfN/8/rStljEqy5PuJUdIWy9zIaMUI+4oSeJWKVACkCyG2VryUqM
D79+4xzf4XqvpH1OLu+jmcWofYougFJdUFv4gFzofMMTgnygpt01bhip1WvXQX4U
W7URmllhisvTy5+7wd2UraBHBxvg92QmW7EYojerK6Mw8ejpWJcz9DCT3ZolhNxC
REd5ak32XSDXYJkvk2V7Dpq7uL8pqAPvgUKmdFckJ6I+TTn+IdDw7xsHK8Bww2We
c3R3ivIbi1MhXBBR2I//jbLX9ex8jhK7vEVT+8B2tWuOY8DVomziW0ksO87bm+WH
flOE3jkr2ITWB6bqwauto4z42svCdIy8DAVbT0vGlXYQAX2uLPLYsBgVeRvJfJGz
tHkPNgn6vLSgxxwPfr44NkZZt7JG8elsGTpuqapKIf8ttnvV6V9VLLx4muFSIKNO
GnNp3ls/JqSLI7nBD4hqFbK0pqiwgzqHP7oNoeuu88awPJAfAhJboO44pfH8gpXR
W33X3DNQKvIU9yhKXlqbFxBRVbZze3HXdpiLq8uuHpewlWxHwEwR0kmI63jwcyNr
f+RobZgMkjvP3lTWYLhssHYJgggvgcX0myEzZT12u0ibn38w2YPQs+zKs9z7okIX
YWas/df+2XnHvIdlXnjD+dksJzoMuCmxYbCgx5pD/p2qOzuRlqqRjLZs2kem5JJ6
JeVBizD7kyyCDYcFkFKjgpogQHSHXSO9rZq7oWlA5zMk/rFNeFM9uCNdObxt1afb
yi93eMxWqFlaw41iGkHCWDtqGtU5jiZAVd0GvN+B2IgTVIsgAnvntIwn135HGmp4
utrcneXvNeSCqwju6hA00Sll0N92Nh5MjN5dI6nFsGryXG+plf29Pw0kEDe1OVZk
VHMEfRGyyJlM+LBSDWmM8C8oBERbJy5dRuBJJmpcCfWhau5JSTqL9iGqLuPV4AGt
xFGPMsaXJB1WEQGyU5uvHmxtbU8kqOnqkXnDn89mrk7DmLDWPUyaUobwVZ2EJ9dy
noQMv/qY4ljnBPt9404uV9Aq3sevJRE5vihv0lCuj0YtzdeXTFHvRzw8aqppZoat
PLSNs8DK34C0x1lJpkQNu6y1sGZIQo6EZrcQ5+Mp4xZ6ofWmENGmt0OKw6GWK9iF
tciGtRVBzh8BxY7QbgGtqaqftjHroj1XD2vO+D5cJmrw7TB7aNjp08ARrtz+yOZE
HFxz740kiqFHrOAJK6Lgi94RecfPQx4gM15kxCh8Bgy0h5NPa5ZscbkxBfTs6TYt
SxowywaI/7RJC2nJ5SDgUIrA085H0N+1IJOlaaiV3+iQef3znaNS7sSagucjj5NI
jJAA3eGexL/dZ6j57iQk5TR7CXcXAVFikv9nX1+hUGyEM5ZmKPo9gO90PklMKyoP
lefy+pB+on0CN7+x+pxx7vbo+OrvuvvMq8FIwgdXWvVmpl1+peK9LNxuSklCg5bf
7s1RJ7VhfLMYmfT+2GxPg8751jgrUWfl5ebuXAI0ROfSOCt96qNTqQ5gMZlFDlaU
NSXtbmuUYp1xwRi455pmdyyvI8BpADeEAcsy2cmaYaJZVBQMQxYkHq8ZVYh3A/6F
RqY8Es7K6OTRHcVbF6HTxQm5gAppfVveHk9KI7s5XSePujBO02LiLTotZmgegBCn
6TglWWmYBVmoYE6J4gm+U/KVPBj8hlQdKbNSg7B3/xmK9zvq6uM+yx0f3yUg2A7K
1nozEY+CD/L9vmnPiGP5uRqZel612RgEHl263CswoAw7URR/hgYGtYBE51gdidFZ
zj3GkwJnnQleMyizwbLa92kNRLJVOddGZbyIJQvXXbwa3JuHwlcPFoxWFRtqLC7I
DxFw+XpIuHRBNfpr3Wcm3vKE5uAjnObZ9NG+ic/9fPX6s/5ZvBd4plYO5FLOwAye
P7+r4R+Zog5RFwSfFnhurJBleg83fRlyjr8pF+uopv1WYBCpMhS8ETTAsRkCvIk9
A411LXSaD5b8P5rEDvOPlW1AHIiKoisbLpXhKQw8hTQwtVJ7A9sr3w9Sj76YW48S
TykaM5SWyfSHeRWkZvFAFM2DQ/HnxQ909QBwW7InKmtmmMcHDfLyNArKsQuFk3j2
6B2coqbf8tmvSf7s6JGPs0HCjHPUPRwiadJepwLqn0n5YscqzKkc0tpgDMhtqLxV
7r3gfT2TPppIsm+iYRlVAUWMBYQNeAcAoqr35B9e6ZagUE0X0zVInid3yVjbg3Pr
JgX2PB8NTaSIScJBcWmX9CYG0f1L8G/C4E9kB9JwZDClFN+ADrLaTwSy0laW2T+2
VLa3y36tY/3x3+o0RP1VBS3SyM1ZLtiwLIDVJBACZmgObu3DpcuGedIvIUvgjTUQ
zXDmGURaqs4LaNdIFpqy0YKCmmmQ1d1n2Gt00u+jQAizBXI0h1pYOf8XRb+u9e67
Yzt81BCRR6dyQ5Bc/FbGjO/9ObT/TI9JhHy5wKBvCVwzV0swrdxw5Z+KqE0NpcXM
r/hHIj5w9kPTrl+49v5b2IWoq0E2LtiCCu8RqeDL3C+I60OIUWsuzdXT+oRAlDaB
5/qmXdcGzyIxiKvafNfcV8x+wVEabx3bDm4jwgE3b2PX5u8vJHcSam/itjISnCfi
thk5CEhUzNV9VQDGy4+MaQP26l/ycz/4E02+IqCL+K5ewsPAgEdDOkpXL6ICTmkk
1YjCc1Dj9iaMk9vuS+0F5v6m9z+vOxn7tXvS/3wm+11x7MnUqqzdtKkCuvS5/nHv
A8dM4jFmT7bn08C6frugv8RX9yXy4KQv/8Y4+57Aj8vomdtqhgF6Q8IhWDi0uFT6
2m8Vxz59K4WkVhvCQM7hhTVGVxfuQwmhXqQE/f0d5X4CLVwaBPaHPu0VdEwQ+hU9
qoMPAC0jmmcJgfRKMxsFpCLmNw7h4//WBzUZeuUsW56lYQ3wvWETC8kzMs834N6q
M67UGmc8uzeDT8wdvptRroB2yVNl4WiWoQUXnsszyud00amsn4gklQDbQAuVKimb
3d36y6RMmbkLMr9HTQ/Qqr6lpi8TAR3+/CK5S3aBEv/cZickxZPazUz9I6vEURJ1
EyRQyr/TYyLSXG5WPc4p9BMon1qGD0VMlsn3G1fA3Fv+e9vx+aMdI3LLto5iOSR6
za3Ld60X+auphGsmIomXs15pTLST1g96YrTShw1ZjL50144TgRAQ68UhmT7lXlvi
JWUpeZZzeZAFbddZagKM82ncNIsLNymWWObwkbvsYZaTSKhKseIppF1I+i4QTv7q
ru7sgMzF7oRpMnezPDLEFnCO+VZS8WWk1FgXYneujZnySKQdpfeDhEk8/Mn7xC5k
4iGaURTz6gKoIsxhpkQIfiQbRhncA2BMXxNhP/Iltmvqq/h9rYxd3L11dE8OWavb
nF9R1kB47Fqary0bt2sw0ksOsN6UOkCmJcwa11+nL3AMOG5sskHWXa7Cm2La2aYM
26Ke5jIBmqW0YyjjB8xw+Xmo1EXrjPbZeLA3qam+/eM+jq2+9EGZ9ZoDWPjTw2ZG
sMS49XRniOpukUY/GWdkJTtHEmIls4uu58ugJKA0ambE9uWdGZCcgdXKezGIT/vg
d8pLw4TRa6hzSj0vyvvs9a/pZ0+xAhDwd1n95M+GQWa59thlhCcX9fEOVbWge+Ag
+C5ypg4M3USEVDuqgNsqB8XPHvUZ9lJT94IQpL0Jk5I6M5QURMBzpCnSH0veUa4q
TZ1pb+kvWj0E1CRfteQTGNjBgJVrR8KaRSQ14nluWrSpGjBPEIfd1mYn+IKETc88
sX6NJZgfC+SmZ0pea7hDqjFtfWfxGZXoaIREH7WHQpIfxWrDb0xKUyfwe0O7UHIg
Vi7zD0/HqEFb484u+Xv9ytKcDVAj8oCvHD0VkJU+aFUxK+mZVRXtEk7UZ1VVh8/i
ndY9er48yLsrTNpprJT33GaMtWcz/Z6UwxMKtz0MYf+bPFAVObzHWC9rxXfsiPUY
7PlQDebBdmAku+kCbFtEZ24TcjrMVpNQel72LMT4sxN6qjCEFFKhSOEpJgO1L1mI
q6lJ/OruOQkQuTwVTk/T8Jk5uc4fXhwB75TIXE9BpcJPEBN0kVYT3REWfFhsaizY
QU+QWW6MpL1ary3gI7NsBGAVxSUPRTQ+90LWclkNqUyeF+HDY5us7ZIAIiexuUDm
BLEOpngRtwLEMr0xWWADP1Kimp9CGf4Np3Pjj0hSFkHICnx8JVDKcg5zLjv8NMyd
SqoZPd/sFj5SBmn6PIK2G91183XXSDttA//5N7bq3dFp9aQs9lVWqTMuMoAraAe+
kVHK4roL5+i4RZ8HSuPIv5gTe9vDgMaHDWIxhK+mJi3znKGy9mOxjWP1DeO4AiXm
vxuRWToknwT+E7KDz/N5m9Sp0HajdJIwLQpq/lJ5amuJ4kKTeJVnoHWVjQ+Rtkqa
tJdcF5OViCCgTZAVHZhJHscu8y22IMTcL4yFtYctlTx+P8vDJ+xtlvOq02nyk4RH
ROOs7knQDh9LykQw4WOqOxmii2lK/b7GtRuMsddgkk6vnHuehlZNaeksow+yw3Px
MVCdMGg9Xd6WMWFiJBQCm1UN5GWqfXTVUOK1m2SVwrG7BoB4dlndjxZXKgtEJEVV
6AM0qDFlzrS8h4BhXNQFSG26Bod8ba8l3bjjiNJfb9wlyW72bgFqxAq+tQD1lZxj
urtrIYLBMir0JupOhswH3LtspdGnOizpq2hg2MGtZ4Mpv+piMdvV6HYsfDF22XwB
3spv0SavpaBBAsQK9En6zKF7XXVlCjiiwa06zD3FRaLo3dWTPHr+Dx7uzreQ/nqR
27R7OVeWhK6DVZfgabql9ouRGkuvsogCfXSwLhQBbpokNFjwQC50LwHNQvMZ62zM
vVC+m1XU7YaHri1QQXyQz2j/x4o+b8hqxwZr9pkcCdO8Wv9RGC5ewqcYRn0Qza/p
+XqKCCIuqebLus/AF6D2/4YGmIJoJJAL3vWXjVDtHl79YpnOacIHjfMDlwfG/Hkk
FC3kRvbidi3tmgwPisAiytWh2guZD72XgUETehLcpmSt/onSHySMwrHO1/k87UuX
`pragma protect end_protected
